module sign_mag_adder_lut #(
    parameter WIDTH = 8
) (
    input  logic             clk,
    input  logic [WIDTH-1:0] a_in,
    input  logic [WIDTH-1:0] b_in,
    output logic [WIDTH-1:0] adder_out
);
    logic [WIDTH-1:0] data_out;

    generate
        if (WIDTH == 4)
        begin
            always_comb 
            begin
                case({a_in, b_in})
                    8'h00: data_out = 4'h0;
                    8'h01: data_out = 4'h1;
                    8'h02: data_out = 4'h2;
                    8'h03: data_out = 4'h3;
                    8'h04: data_out = 4'h4;
                    8'h05: data_out = 4'h5;
                    8'h06: data_out = 4'h6;
                    8'h07: data_out = 4'h7;
                    8'h08: data_out = 4'h0;
                    8'h09: data_out = 4'h9;
                    8'h0A: data_out = 4'hA;
                    8'h0B: data_out = 4'hB;
                    8'h0C: data_out = 4'hC;
                    8'h0D: data_out = 4'hD;
                    8'h0E: data_out = 4'hE;
                    8'h0F: data_out = 4'hF;
                    8'h10: data_out = 4'h1;
                    8'h11: data_out = 4'h2;
                    8'h12: data_out = 4'h3;
                    8'h13: data_out = 4'h4;
                    8'h14: data_out = 4'h5;
                    8'h15: data_out = 4'h6;
                    8'h16: data_out = 4'h7;
                    8'h17: data_out = 4'h8;
                    8'h18: data_out = 4'h1;
                    8'h19: data_out = 4'h0;
                    8'h1A: data_out = 4'h9;
                    8'h1B: data_out = 4'hA;
                    8'h1C: data_out = 4'hB;
                    8'h1D: data_out = 4'hC;
                    8'h1E: data_out = 4'hD;
                    8'h1F: data_out = 4'hE;
                    8'h20: data_out = 4'h2;
                    8'h21: data_out = 4'h3;
                    8'h22: data_out = 4'h4;
                    8'h23: data_out = 4'h5;
                    8'h24: data_out = 4'h6;
                    8'h25: data_out = 4'h7;
                    8'h26: data_out = 4'h8;
                    8'h27: data_out = 4'h9;
                    8'h28: data_out = 4'h2;
                    8'h29: data_out = 4'h1;
                    8'h2A: data_out = 4'h0;
                    8'h2B: data_out = 4'h9;
                    8'h2C: data_out = 4'hA;
                    8'h2D: data_out = 4'hB;
                    8'h2E: data_out = 4'hC;
                    8'h2F: data_out = 4'hD;
                    8'h30: data_out = 4'h3;
                    8'h31: data_out = 4'h4;
                    8'h32: data_out = 4'h5;
                    8'h33: data_out = 4'h6;
                    8'h34: data_out = 4'h7;
                    8'h35: data_out = 4'h8;
                    8'h36: data_out = 4'h9;
                    8'h37: data_out = 4'hA;
                    8'h38: data_out = 4'h3;
                    8'h39: data_out = 4'h2;
                    8'h3A: data_out = 4'h1;
                    8'h3B: data_out = 4'h0;
                    8'h3C: data_out = 4'h9;
                    8'h3D: data_out = 4'hA;
                    8'h3E: data_out = 4'hB;
                    8'h3F: data_out = 4'hC;
                    8'h40: data_out = 4'h4;
                    8'h41: data_out = 4'h5;
                    8'h42: data_out = 4'h6;
                    8'h43: data_out = 4'h7;
                    8'h44: data_out = 4'h8;
                    8'h45: data_out = 4'h9;
                    8'h46: data_out = 4'hA;
                    8'h47: data_out = 4'hB;
                    8'h48: data_out = 4'h4;
                    8'h49: data_out = 4'h3;
                    8'h4A: data_out = 4'h2;
                    8'h4B: data_out = 4'h1;
                    8'h4C: data_out = 4'h0;
                    8'h4D: data_out = 4'h9;
                    8'h4E: data_out = 4'hA;
                    8'h4F: data_out = 4'hB;
                    8'h50: data_out = 4'h5;
                    8'h51: data_out = 4'h6;
                    8'h52: data_out = 4'h7;
                    8'h53: data_out = 4'h8;
                    8'h54: data_out = 4'h9;
                    8'h55: data_out = 4'hA;
                    8'h56: data_out = 4'hB;
                    8'h57: data_out = 4'hC;
                    8'h58: data_out = 4'h5;
                    8'h59: data_out = 4'h4;
                    8'h5A: data_out = 4'h3;
                    8'h5B: data_out = 4'h2;
                    8'h5C: data_out = 4'h1;
                    8'h5D: data_out = 4'h0;
                    8'h5E: data_out = 4'h9;
                    8'h5F: data_out = 4'hA;
                    8'h60: data_out = 4'h6;
                    8'h61: data_out = 4'h7;
                    8'h62: data_out = 4'h8;
                    8'h63: data_out = 4'h9;
                    8'h64: data_out = 4'hA;
                    8'h65: data_out = 4'hB;
                    8'h66: data_out = 4'hC;
                    8'h67: data_out = 4'hD;
                    8'h68: data_out = 4'h6;
                    8'h69: data_out = 4'h5;
                    8'h6A: data_out = 4'h4;
                    8'h6B: data_out = 4'h3;
                    8'h6C: data_out = 4'h2;
                    8'h6D: data_out = 4'h1;
                    8'h6E: data_out = 4'h0;
                    8'h6F: data_out = 4'h9;
                    8'h70: data_out = 4'h7;
                    8'h71: data_out = 4'h8;
                    8'h72: data_out = 4'h9;
                    8'h73: data_out = 4'hA;
                    8'h74: data_out = 4'hB;
                    8'h75: data_out = 4'hC;
                    8'h76: data_out = 4'hD;
                    8'h77: data_out = 4'hE;
                    8'h78: data_out = 4'h7;
                    8'h79: data_out = 4'h6;
                    8'h7A: data_out = 4'h5;
                    8'h7B: data_out = 4'h4;
                    8'h7C: data_out = 4'h3;
                    8'h7D: data_out = 4'h2;
                    8'h7E: data_out = 4'h1;
                    8'h7F: data_out = 4'h0;
                    8'h80: data_out = 4'h0;
                    8'h81: data_out = 4'h1;
                    8'h82: data_out = 4'h2;
                    8'h83: data_out = 4'h3;
                    8'h84: data_out = 4'h4;
                    8'h85: data_out = 4'h5;
                    8'h86: data_out = 4'h6;
                    8'h87: data_out = 4'h7;
                    8'h88: data_out = 4'h0;
                    8'h89: data_out = 4'h9;
                    8'h8A: data_out = 4'hA;
                    8'h8B: data_out = 4'hB;
                    8'h8C: data_out = 4'hC;
                    8'h8D: data_out = 4'hD;
                    8'h8E: data_out = 4'hE;
                    8'h8F: data_out = 4'hF;
                    8'h90: data_out = 4'h9;
                    8'h91: data_out = 4'h0;
                    8'h92: data_out = 4'h1;
                    8'h93: data_out = 4'h2;
                    8'h94: data_out = 4'h3;
                    8'h95: data_out = 4'h4;
                    8'h96: data_out = 4'h5;
                    8'h97: data_out = 4'h6;
                    8'h98: data_out = 4'h9;
                    8'h99: data_out = 4'hA;
                    8'h9A: data_out = 4'hB;
                    8'h9B: data_out = 4'hC;
                    8'h9C: data_out = 4'hD;
                    8'h9D: data_out = 4'hE;
                    8'h9E: data_out = 4'hF;
                    8'h9F: data_out = 4'h8;
                    8'hA0: data_out = 4'hA;
                    8'hA1: data_out = 4'h9;
                    8'hA2: data_out = 4'h0;
                    8'hA3: data_out = 4'h1;
                    8'hA4: data_out = 4'h2;
                    8'hA5: data_out = 4'h3;
                    8'hA6: data_out = 4'h4;
                    8'hA7: data_out = 4'h5;
                    8'hA8: data_out = 4'hA;
                    8'hA9: data_out = 4'hB;
                    8'hAA: data_out = 4'hC;
                    8'hAB: data_out = 4'hD;
                    8'hAC: data_out = 4'hE;
                    8'hAD: data_out = 4'hF;
                    8'hAE: data_out = 4'h8;
                    8'hAF: data_out = 4'h9;
                    8'hB0: data_out = 4'hB;
                    8'hB1: data_out = 4'hA;
                    8'hB2: data_out = 4'h9;
                    8'hB3: data_out = 4'h0;
                    8'hB4: data_out = 4'h1;
                    8'hB5: data_out = 4'h2;
                    8'hB6: data_out = 4'h3;
                    8'hB7: data_out = 4'h4;
                    8'hB8: data_out = 4'hB;
                    8'hB9: data_out = 4'hC;
                    8'hBA: data_out = 4'hD;
                    8'hBB: data_out = 4'hE;
                    8'hBC: data_out = 4'hF;
                    8'hBD: data_out = 4'h8;
                    8'hBE: data_out = 4'h9;
                    8'hBF: data_out = 4'hA;
                    8'hC0: data_out = 4'hC;
                    8'hC1: data_out = 4'hB;
                    8'hC2: data_out = 4'hA;
                    8'hC3: data_out = 4'h9;
                    8'hC4: data_out = 4'h0;
                    8'hC5: data_out = 4'h1;
                    8'hC6: data_out = 4'h2;
                    8'hC7: data_out = 4'h3;
                    8'hC8: data_out = 4'hC;
                    8'hC9: data_out = 4'hD;
                    8'hCA: data_out = 4'hE;
                    8'hCB: data_out = 4'hF;
                    8'hCC: data_out = 4'h8;
                    8'hCD: data_out = 4'h9;
                    8'hCE: data_out = 4'hA;
                    8'hCF: data_out = 4'hB;
                    8'hD0: data_out = 4'hD;
                    8'hD1: data_out = 4'hC;
                    8'hD2: data_out = 4'hB;
                    8'hD3: data_out = 4'hA;
                    8'hD4: data_out = 4'h9;
                    8'hD5: data_out = 4'h0;
                    8'hD6: data_out = 4'h1;
                    8'hD7: data_out = 4'h2;
                    8'hD8: data_out = 4'hD;
                    8'hD9: data_out = 4'hE;
                    8'hDA: data_out = 4'hF;
                    8'hDB: data_out = 4'h8;
                    8'hDC: data_out = 4'h9;
                    8'hDD: data_out = 4'hA;
                    8'hDE: data_out = 4'hB;
                    8'hDF: data_out = 4'hC;
                    8'hE0: data_out = 4'hE;
                    8'hE1: data_out = 4'hD;
                    8'hE2: data_out = 4'hC;
                    8'hE3: data_out = 4'hB;
                    8'hE4: data_out = 4'hA;
                    8'hE5: data_out = 4'h9;
                    8'hE6: data_out = 4'h0;
                    8'hE7: data_out = 4'h1;
                    8'hE8: data_out = 4'hE;
                    8'hE9: data_out = 4'hF;
                    8'hEA: data_out = 4'h8;
                    8'hEB: data_out = 4'h9;
                    8'hEC: data_out = 4'hA;
                    8'hED: data_out = 4'hB;
                    8'hEE: data_out = 4'hC;
                    8'hEF: data_out = 4'hD;
                    8'hF0: data_out = 4'hF;
                    8'hF1: data_out = 4'hE;
                    8'hF2: data_out = 4'hD;
                    8'hF3: data_out = 4'hC;
                    8'hF4: data_out = 4'hB;
                    8'hF5: data_out = 4'hA;
                    8'hF6: data_out = 4'h9;
                    8'hF7: data_out = 4'h0;
                    8'hF8: data_out = 4'hF;
                    8'hF9: data_out = 4'h8;
                    8'hFA: data_out = 4'h9;
                    8'hFB: data_out = 4'hA;
                    8'hFC: data_out = 4'hB;
                    8'hFD: data_out = 4'hC;
                    8'hFE: data_out = 4'hD;
                    8'hFF: data_out = 4'hE;
                    default: data_out = 4'h0;
                endcase
            end
        end
        else
        begin
            always_comb 
            begin : ROM_blk
                case({a_in, b_in})
                    16'h0000: data_out = 8'h0;
                    16'h0001: data_out = 8'h1;
                    16'h0002: data_out = 8'h2;
                    16'h0003: data_out = 8'h3;
                    16'h0004: data_out = 8'h4;
                    16'h0005: data_out = 8'h5;
                    16'h0006: data_out = 8'h6;
                    16'h0007: data_out = 8'h7;
                    16'h0008: data_out = 8'h8;
                    16'h0009: data_out = 8'h9;
                    16'h000A: data_out = 8'hA;
                    16'h000B: data_out = 8'hB;
                    16'h000C: data_out = 8'hC;
                    16'h000D: data_out = 8'hD;
                    16'h000E: data_out = 8'hE;
                    16'h000F: data_out = 8'hF;
                    16'h0010: data_out = 8'h10;
                    16'h0011: data_out = 8'h11;
                    16'h0012: data_out = 8'h12;
                    16'h0013: data_out = 8'h13;
                    16'h0014: data_out = 8'h14;
                    16'h0015: data_out = 8'h15;
                    16'h0016: data_out = 8'h16;
                    16'h0017: data_out = 8'h17;
                    16'h0018: data_out = 8'h18;
                    16'h0019: data_out = 8'h19;
                    16'h001A: data_out = 8'h1A;
                    16'h001B: data_out = 8'h1B;
                    16'h001C: data_out = 8'h1C;
                    16'h001D: data_out = 8'h1D;
                    16'h001E: data_out = 8'h1E;
                    16'h001F: data_out = 8'h1F;
                    16'h0020: data_out = 8'h20;
                    16'h0021: data_out = 8'h21;
                    16'h0022: data_out = 8'h22;
                    16'h0023: data_out = 8'h23;
                    16'h0024: data_out = 8'h24;
                    16'h0025: data_out = 8'h25;
                    16'h0026: data_out = 8'h26;
                    16'h0027: data_out = 8'h27;
                    16'h0028: data_out = 8'h28;
                    16'h0029: data_out = 8'h29;
                    16'h002A: data_out = 8'h2A;
                    16'h002B: data_out = 8'h2B;
                    16'h002C: data_out = 8'h2C;
                    16'h002D: data_out = 8'h2D;
                    16'h002E: data_out = 8'h2E;
                    16'h002F: data_out = 8'h2F;
                    16'h0030: data_out = 8'h30;
                    16'h0031: data_out = 8'h31;
                    16'h0032: data_out = 8'h32;
                    16'h0033: data_out = 8'h33;
                    16'h0034: data_out = 8'h34;
                    16'h0035: data_out = 8'h35;
                    16'h0036: data_out = 8'h36;
                    16'h0037: data_out = 8'h37;
                    16'h0038: data_out = 8'h38;
                    16'h0039: data_out = 8'h39;
                    16'h003A: data_out = 8'h3A;
                    16'h003B: data_out = 8'h3B;
                    16'h003C: data_out = 8'h3C;
                    16'h003D: data_out = 8'h3D;
                    16'h003E: data_out = 8'h3E;
                    16'h003F: data_out = 8'h3F;
                    16'h0040: data_out = 8'h40;
                    16'h0041: data_out = 8'h41;
                    16'h0042: data_out = 8'h42;
                    16'h0043: data_out = 8'h43;
                    16'h0044: data_out = 8'h44;
                    16'h0045: data_out = 8'h45;
                    16'h0046: data_out = 8'h46;
                    16'h0047: data_out = 8'h47;
                    16'h0048: data_out = 8'h48;
                    16'h0049: data_out = 8'h49;
                    16'h004A: data_out = 8'h4A;
                    16'h004B: data_out = 8'h4B;
                    16'h004C: data_out = 8'h4C;
                    16'h004D: data_out = 8'h4D;
                    16'h004E: data_out = 8'h4E;
                    16'h004F: data_out = 8'h4F;
                    16'h0050: data_out = 8'h50;
                    16'h0051: data_out = 8'h51;
                    16'h0052: data_out = 8'h52;
                    16'h0053: data_out = 8'h53;
                    16'h0054: data_out = 8'h54;
                    16'h0055: data_out = 8'h55;
                    16'h0056: data_out = 8'h56;
                    16'h0057: data_out = 8'h57;
                    16'h0058: data_out = 8'h58;
                    16'h0059: data_out = 8'h59;
                    16'h005A: data_out = 8'h5A;
                    16'h005B: data_out = 8'h5B;
                    16'h005C: data_out = 8'h5C;
                    16'h005D: data_out = 8'h5D;
                    16'h005E: data_out = 8'h5E;
                    16'h005F: data_out = 8'h5F;
                    16'h0060: data_out = 8'h60;
                    16'h0061: data_out = 8'h61;
                    16'h0062: data_out = 8'h62;
                    16'h0063: data_out = 8'h63;
                    16'h0064: data_out = 8'h64;
                    16'h0065: data_out = 8'h65;
                    16'h0066: data_out = 8'h66;
                    16'h0067: data_out = 8'h67;
                    16'h0068: data_out = 8'h68;
                    16'h0069: data_out = 8'h69;
                    16'h006A: data_out = 8'h6A;
                    16'h006B: data_out = 8'h6B;
                    16'h006C: data_out = 8'h6C;
                    16'h006D: data_out = 8'h6D;
                    16'h006E: data_out = 8'h6E;
                    16'h006F: data_out = 8'h6F;
                    16'h0070: data_out = 8'h70;
                    16'h0071: data_out = 8'h71;
                    16'h0072: data_out = 8'h72;
                    16'h0073: data_out = 8'h73;
                    16'h0074: data_out = 8'h74;
                    16'h0075: data_out = 8'h75;
                    16'h0076: data_out = 8'h76;
                    16'h0077: data_out = 8'h77;
                    16'h0078: data_out = 8'h78;
                    16'h0079: data_out = 8'h79;
                    16'h007A: data_out = 8'h7A;
                    16'h007B: data_out = 8'h7B;
                    16'h007C: data_out = 8'h7C;
                    16'h007D: data_out = 8'h7D;
                    16'h007E: data_out = 8'h7E;
                    16'h007F: data_out = 8'h7F;
                    16'h0080: data_out = 8'h0;
                    16'h0081: data_out = 8'h81;
                    16'h0082: data_out = 8'h82;
                    16'h0083: data_out = 8'h83;
                    16'h0084: data_out = 8'h84;
                    16'h0085: data_out = 8'h85;
                    16'h0086: data_out = 8'h86;
                    16'h0087: data_out = 8'h87;
                    16'h0088: data_out = 8'h88;
                    16'h0089: data_out = 8'h89;
                    16'h008A: data_out = 8'h8A;
                    16'h008B: data_out = 8'h8B;
                    16'h008C: data_out = 8'h8C;
                    16'h008D: data_out = 8'h8D;
                    16'h008E: data_out = 8'h8E;
                    16'h008F: data_out = 8'h8F;
                    16'h0090: data_out = 8'h90;
                    16'h0091: data_out = 8'h91;
                    16'h0092: data_out = 8'h92;
                    16'h0093: data_out = 8'h93;
                    16'h0094: data_out = 8'h94;
                    16'h0095: data_out = 8'h95;
                    16'h0096: data_out = 8'h96;
                    16'h0097: data_out = 8'h97;
                    16'h0098: data_out = 8'h98;
                    16'h0099: data_out = 8'h99;
                    16'h009A: data_out = 8'h9A;
                    16'h009B: data_out = 8'h9B;
                    16'h009C: data_out = 8'h9C;
                    16'h009D: data_out = 8'h9D;
                    16'h009E: data_out = 8'h9E;
                    16'h009F: data_out = 8'h9F;
                    16'h00A0: data_out = 8'hA0;
                    16'h00A1: data_out = 8'hA1;
                    16'h00A2: data_out = 8'hA2;
                    16'h00A3: data_out = 8'hA3;
                    16'h00A4: data_out = 8'hA4;
                    16'h00A5: data_out = 8'hA5;
                    16'h00A6: data_out = 8'hA6;
                    16'h00A7: data_out = 8'hA7;
                    16'h00A8: data_out = 8'hA8;
                    16'h00A9: data_out = 8'hA9;
                    16'h00AA: data_out = 8'hAA;
                    16'h00AB: data_out = 8'hAB;
                    16'h00AC: data_out = 8'hAC;
                    16'h00AD: data_out = 8'hAD;
                    16'h00AE: data_out = 8'hAE;
                    16'h00AF: data_out = 8'hAF;
                    16'h00B0: data_out = 8'hB0;
                    16'h00B1: data_out = 8'hB1;
                    16'h00B2: data_out = 8'hB2;
                    16'h00B3: data_out = 8'hB3;
                    16'h00B4: data_out = 8'hB4;
                    16'h00B5: data_out = 8'hB5;
                    16'h00B6: data_out = 8'hB6;
                    16'h00B7: data_out = 8'hB7;
                    16'h00B8: data_out = 8'hB8;
                    16'h00B9: data_out = 8'hB9;
                    16'h00BA: data_out = 8'hBA;
                    16'h00BB: data_out = 8'hBB;
                    16'h00BC: data_out = 8'hBC;
                    16'h00BD: data_out = 8'hBD;
                    16'h00BE: data_out = 8'hBE;
                    16'h00BF: data_out = 8'hBF;
                    16'h00C0: data_out = 8'hC0;
                    16'h00C1: data_out = 8'hC1;
                    16'h00C2: data_out = 8'hC2;
                    16'h00C3: data_out = 8'hC3;
                    16'h00C4: data_out = 8'hC4;
                    16'h00C5: data_out = 8'hC5;
                    16'h00C6: data_out = 8'hC6;
                    16'h00C7: data_out = 8'hC7;
                    16'h00C8: data_out = 8'hC8;
                    16'h00C9: data_out = 8'hC9;
                    16'h00CA: data_out = 8'hCA;
                    16'h00CB: data_out = 8'hCB;
                    16'h00CC: data_out = 8'hCC;
                    16'h00CD: data_out = 8'hCD;
                    16'h00CE: data_out = 8'hCE;
                    16'h00CF: data_out = 8'hCF;
                    16'h00D0: data_out = 8'hD0;
                    16'h00D1: data_out = 8'hD1;
                    16'h00D2: data_out = 8'hD2;
                    16'h00D3: data_out = 8'hD3;
                    16'h00D4: data_out = 8'hD4;
                    16'h00D5: data_out = 8'hD5;
                    16'h00D6: data_out = 8'hD6;
                    16'h00D7: data_out = 8'hD7;
                    16'h00D8: data_out = 8'hD8;
                    16'h00D9: data_out = 8'hD9;
                    16'h00DA: data_out = 8'hDA;
                    16'h00DB: data_out = 8'hDB;
                    16'h00DC: data_out = 8'hDC;
                    16'h00DD: data_out = 8'hDD;
                    16'h00DE: data_out = 8'hDE;
                    16'h00DF: data_out = 8'hDF;
                    16'h00E0: data_out = 8'hE0;
                    16'h00E1: data_out = 8'hE1;
                    16'h00E2: data_out = 8'hE2;
                    16'h00E3: data_out = 8'hE3;
                    16'h00E4: data_out = 8'hE4;
                    16'h00E5: data_out = 8'hE5;
                    16'h00E6: data_out = 8'hE6;
                    16'h00E7: data_out = 8'hE7;
                    16'h00E8: data_out = 8'hE8;
                    16'h00E9: data_out = 8'hE9;
                    16'h00EA: data_out = 8'hEA;
                    16'h00EB: data_out = 8'hEB;
                    16'h00EC: data_out = 8'hEC;
                    16'h00ED: data_out = 8'hED;
                    16'h00EE: data_out = 8'hEE;
                    16'h00EF: data_out = 8'hEF;
                    16'h00F0: data_out = 8'hF0;
                    16'h00F1: data_out = 8'hF1;
                    16'h00F2: data_out = 8'hF2;
                    16'h00F3: data_out = 8'hF3;
                    16'h00F4: data_out = 8'hF4;
                    16'h00F5: data_out = 8'hF5;
                    16'h00F6: data_out = 8'hF6;
                    16'h00F7: data_out = 8'hF7;
                    16'h00F8: data_out = 8'hF8;
                    16'h00F9: data_out = 8'hF9;
                    16'h00FA: data_out = 8'hFA;
                    16'h00FB: data_out = 8'hFB;
                    16'h00FC: data_out = 8'hFC;
                    16'h00FD: data_out = 8'hFD;
                    16'h00FE: data_out = 8'hFE;
                    16'h00FF: data_out = 8'hFF;
                    16'h0100: data_out = 8'h1;
                    16'h0101: data_out = 8'h2;
                    16'h0102: data_out = 8'h3;
                    16'h0103: data_out = 8'h4;
                    16'h0104: data_out = 8'h5;
                    16'h0105: data_out = 8'h6;
                    16'h0106: data_out = 8'h7;
                    16'h0107: data_out = 8'h8;
                    16'h0108: data_out = 8'h9;
                    16'h0109: data_out = 8'hA;
                    16'h010A: data_out = 8'hB;
                    16'h010B: data_out = 8'hC;
                    16'h010C: data_out = 8'hD;
                    16'h010D: data_out = 8'hE;
                    16'h010E: data_out = 8'hF;
                    16'h010F: data_out = 8'h10;
                    16'h0110: data_out = 8'h11;
                    16'h0111: data_out = 8'h12;
                    16'h0112: data_out = 8'h13;
                    16'h0113: data_out = 8'h14;
                    16'h0114: data_out = 8'h15;
                    16'h0115: data_out = 8'h16;
                    16'h0116: data_out = 8'h17;
                    16'h0117: data_out = 8'h18;
                    16'h0118: data_out = 8'h19;
                    16'h0119: data_out = 8'h1A;
                    16'h011A: data_out = 8'h1B;
                    16'h011B: data_out = 8'h1C;
                    16'h011C: data_out = 8'h1D;
                    16'h011D: data_out = 8'h1E;
                    16'h011E: data_out = 8'h1F;
                    16'h011F: data_out = 8'h20;
                    16'h0120: data_out = 8'h21;
                    16'h0121: data_out = 8'h22;
                    16'h0122: data_out = 8'h23;
                    16'h0123: data_out = 8'h24;
                    16'h0124: data_out = 8'h25;
                    16'h0125: data_out = 8'h26;
                    16'h0126: data_out = 8'h27;
                    16'h0127: data_out = 8'h28;
                    16'h0128: data_out = 8'h29;
                    16'h0129: data_out = 8'h2A;
                    16'h012A: data_out = 8'h2B;
                    16'h012B: data_out = 8'h2C;
                    16'h012C: data_out = 8'h2D;
                    16'h012D: data_out = 8'h2E;
                    16'h012E: data_out = 8'h2F;
                    16'h012F: data_out = 8'h30;
                    16'h0130: data_out = 8'h31;
                    16'h0131: data_out = 8'h32;
                    16'h0132: data_out = 8'h33;
                    16'h0133: data_out = 8'h34;
                    16'h0134: data_out = 8'h35;
                    16'h0135: data_out = 8'h36;
                    16'h0136: data_out = 8'h37;
                    16'h0137: data_out = 8'h38;
                    16'h0138: data_out = 8'h39;
                    16'h0139: data_out = 8'h3A;
                    16'h013A: data_out = 8'h3B;
                    16'h013B: data_out = 8'h3C;
                    16'h013C: data_out = 8'h3D;
                    16'h013D: data_out = 8'h3E;
                    16'h013E: data_out = 8'h3F;
                    16'h013F: data_out = 8'h40;
                    16'h0140: data_out = 8'h41;
                    16'h0141: data_out = 8'h42;
                    16'h0142: data_out = 8'h43;
                    16'h0143: data_out = 8'h44;
                    16'h0144: data_out = 8'h45;
                    16'h0145: data_out = 8'h46;
                    16'h0146: data_out = 8'h47;
                    16'h0147: data_out = 8'h48;
                    16'h0148: data_out = 8'h49;
                    16'h0149: data_out = 8'h4A;
                    16'h014A: data_out = 8'h4B;
                    16'h014B: data_out = 8'h4C;
                    16'h014C: data_out = 8'h4D;
                    16'h014D: data_out = 8'h4E;
                    16'h014E: data_out = 8'h4F;
                    16'h014F: data_out = 8'h50;
                    16'h0150: data_out = 8'h51;
                    16'h0151: data_out = 8'h52;
                    16'h0152: data_out = 8'h53;
                    16'h0153: data_out = 8'h54;
                    16'h0154: data_out = 8'h55;
                    16'h0155: data_out = 8'h56;
                    16'h0156: data_out = 8'h57;
                    16'h0157: data_out = 8'h58;
                    16'h0158: data_out = 8'h59;
                    16'h0159: data_out = 8'h5A;
                    16'h015A: data_out = 8'h5B;
                    16'h015B: data_out = 8'h5C;
                    16'h015C: data_out = 8'h5D;
                    16'h015D: data_out = 8'h5E;
                    16'h015E: data_out = 8'h5F;
                    16'h015F: data_out = 8'h60;
                    16'h0160: data_out = 8'h61;
                    16'h0161: data_out = 8'h62;
                    16'h0162: data_out = 8'h63;
                    16'h0163: data_out = 8'h64;
                    16'h0164: data_out = 8'h65;
                    16'h0165: data_out = 8'h66;
                    16'h0166: data_out = 8'h67;
                    16'h0167: data_out = 8'h68;
                    16'h0168: data_out = 8'h69;
                    16'h0169: data_out = 8'h6A;
                    16'h016A: data_out = 8'h6B;
                    16'h016B: data_out = 8'h6C;
                    16'h016C: data_out = 8'h6D;
                    16'h016D: data_out = 8'h6E;
                    16'h016E: data_out = 8'h6F;
                    16'h016F: data_out = 8'h70;
                    16'h0170: data_out = 8'h71;
                    16'h0171: data_out = 8'h72;
                    16'h0172: data_out = 8'h73;
                    16'h0173: data_out = 8'h74;
                    16'h0174: data_out = 8'h75;
                    16'h0175: data_out = 8'h76;
                    16'h0176: data_out = 8'h77;
                    16'h0177: data_out = 8'h78;
                    16'h0178: data_out = 8'h79;
                    16'h0179: data_out = 8'h7A;
                    16'h017A: data_out = 8'h7B;
                    16'h017B: data_out = 8'h7C;
                    16'h017C: data_out = 8'h7D;
                    16'h017D: data_out = 8'h7E;
                    16'h017E: data_out = 8'h7F;
                    16'h017F: data_out = 8'h80;
                    16'h0180: data_out = 8'h1;
                    16'h0181: data_out = 8'h0;
                    16'h0182: data_out = 8'h81;
                    16'h0183: data_out = 8'h82;
                    16'h0184: data_out = 8'h83;
                    16'h0185: data_out = 8'h84;
                    16'h0186: data_out = 8'h85;
                    16'h0187: data_out = 8'h86;
                    16'h0188: data_out = 8'h87;
                    16'h0189: data_out = 8'h88;
                    16'h018A: data_out = 8'h89;
                    16'h018B: data_out = 8'h8A;
                    16'h018C: data_out = 8'h8B;
                    16'h018D: data_out = 8'h8C;
                    16'h018E: data_out = 8'h8D;
                    16'h018F: data_out = 8'h8E;
                    16'h0190: data_out = 8'h8F;
                    16'h0191: data_out = 8'h90;
                    16'h0192: data_out = 8'h91;
                    16'h0193: data_out = 8'h92;
                    16'h0194: data_out = 8'h93;
                    16'h0195: data_out = 8'h94;
                    16'h0196: data_out = 8'h95;
                    16'h0197: data_out = 8'h96;
                    16'h0198: data_out = 8'h97;
                    16'h0199: data_out = 8'h98;
                    16'h019A: data_out = 8'h99;
                    16'h019B: data_out = 8'h9A;
                    16'h019C: data_out = 8'h9B;
                    16'h019D: data_out = 8'h9C;
                    16'h019E: data_out = 8'h9D;
                    16'h019F: data_out = 8'h9E;
                    16'h01A0: data_out = 8'h9F;
                    16'h01A1: data_out = 8'hA0;
                    16'h01A2: data_out = 8'hA1;
                    16'h01A3: data_out = 8'hA2;
                    16'h01A4: data_out = 8'hA3;
                    16'h01A5: data_out = 8'hA4;
                    16'h01A6: data_out = 8'hA5;
                    16'h01A7: data_out = 8'hA6;
                    16'h01A8: data_out = 8'hA7;
                    16'h01A9: data_out = 8'hA8;
                    16'h01AA: data_out = 8'hA9;
                    16'h01AB: data_out = 8'hAA;
                    16'h01AC: data_out = 8'hAB;
                    16'h01AD: data_out = 8'hAC;
                    16'h01AE: data_out = 8'hAD;
                    16'h01AF: data_out = 8'hAE;
                    16'h01B0: data_out = 8'hAF;
                    16'h01B1: data_out = 8'hB0;
                    16'h01B2: data_out = 8'hB1;
                    16'h01B3: data_out = 8'hB2;
                    16'h01B4: data_out = 8'hB3;
                    16'h01B5: data_out = 8'hB4;
                    16'h01B6: data_out = 8'hB5;
                    16'h01B7: data_out = 8'hB6;
                    16'h01B8: data_out = 8'hB7;
                    16'h01B9: data_out = 8'hB8;
                    16'h01BA: data_out = 8'hB9;
                    16'h01BB: data_out = 8'hBA;
                    16'h01BC: data_out = 8'hBB;
                    16'h01BD: data_out = 8'hBC;
                    16'h01BE: data_out = 8'hBD;
                    16'h01BF: data_out = 8'hBE;
                    16'h01C0: data_out = 8'hBF;
                    16'h01C1: data_out = 8'hC0;
                    16'h01C2: data_out = 8'hC1;
                    16'h01C3: data_out = 8'hC2;
                    16'h01C4: data_out = 8'hC3;
                    16'h01C5: data_out = 8'hC4;
                    16'h01C6: data_out = 8'hC5;
                    16'h01C7: data_out = 8'hC6;
                    16'h01C8: data_out = 8'hC7;
                    16'h01C9: data_out = 8'hC8;
                    16'h01CA: data_out = 8'hC9;
                    16'h01CB: data_out = 8'hCA;
                    16'h01CC: data_out = 8'hCB;
                    16'h01CD: data_out = 8'hCC;
                    16'h01CE: data_out = 8'hCD;
                    16'h01CF: data_out = 8'hCE;
                    16'h01D0: data_out = 8'hCF;
                    16'h01D1: data_out = 8'hD0;
                    16'h01D2: data_out = 8'hD1;
                    16'h01D3: data_out = 8'hD2;
                    16'h01D4: data_out = 8'hD3;
                    16'h01D5: data_out = 8'hD4;
                    16'h01D6: data_out = 8'hD5;
                    16'h01D7: data_out = 8'hD6;
                    16'h01D8: data_out = 8'hD7;
                    16'h01D9: data_out = 8'hD8;
                    16'h01DA: data_out = 8'hD9;
                    16'h01DB: data_out = 8'hDA;
                    16'h01DC: data_out = 8'hDB;
                    16'h01DD: data_out = 8'hDC;
                    16'h01DE: data_out = 8'hDD;
                    16'h01DF: data_out = 8'hDE;
                    16'h01E0: data_out = 8'hDF;
                    16'h01E1: data_out = 8'hE0;
                    16'h01E2: data_out = 8'hE1;
                    16'h01E3: data_out = 8'hE2;
                    16'h01E4: data_out = 8'hE3;
                    16'h01E5: data_out = 8'hE4;
                    16'h01E6: data_out = 8'hE5;
                    16'h01E7: data_out = 8'hE6;
                    16'h01E8: data_out = 8'hE7;
                    16'h01E9: data_out = 8'hE8;
                    16'h01EA: data_out = 8'hE9;
                    16'h01EB: data_out = 8'hEA;
                    16'h01EC: data_out = 8'hEB;
                    16'h01ED: data_out = 8'hEC;
                    16'h01EE: data_out = 8'hED;
                    16'h01EF: data_out = 8'hEE;
                    16'h01F0: data_out = 8'hEF;
                    16'h01F1: data_out = 8'hF0;
                    16'h01F2: data_out = 8'hF1;
                    16'h01F3: data_out = 8'hF2;
                    16'h01F4: data_out = 8'hF3;
                    16'h01F5: data_out = 8'hF4;
                    16'h01F6: data_out = 8'hF5;
                    16'h01F7: data_out = 8'hF6;
                    16'h01F8: data_out = 8'hF7;
                    16'h01F9: data_out = 8'hF8;
                    16'h01FA: data_out = 8'hF9;
                    16'h01FB: data_out = 8'hFA;
                    16'h01FC: data_out = 8'hFB;
                    16'h01FD: data_out = 8'hFC;
                    16'h01FE: data_out = 8'hFD;
                    16'h01FF: data_out = 8'hFE;
                    16'h0200: data_out = 8'h2;
                    16'h0201: data_out = 8'h3;
                    16'h0202: data_out = 8'h4;
                    16'h0203: data_out = 8'h5;
                    16'h0204: data_out = 8'h6;
                    16'h0205: data_out = 8'h7;
                    16'h0206: data_out = 8'h8;
                    16'h0207: data_out = 8'h9;
                    16'h0208: data_out = 8'hA;
                    16'h0209: data_out = 8'hB;
                    16'h020A: data_out = 8'hC;
                    16'h020B: data_out = 8'hD;
                    16'h020C: data_out = 8'hE;
                    16'h020D: data_out = 8'hF;
                    16'h020E: data_out = 8'h10;
                    16'h020F: data_out = 8'h11;
                    16'h0210: data_out = 8'h12;
                    16'h0211: data_out = 8'h13;
                    16'h0212: data_out = 8'h14;
                    16'h0213: data_out = 8'h15;
                    16'h0214: data_out = 8'h16;
                    16'h0215: data_out = 8'h17;
                    16'h0216: data_out = 8'h18;
                    16'h0217: data_out = 8'h19;
                    16'h0218: data_out = 8'h1A;
                    16'h0219: data_out = 8'h1B;
                    16'h021A: data_out = 8'h1C;
                    16'h021B: data_out = 8'h1D;
                    16'h021C: data_out = 8'h1E;
                    16'h021D: data_out = 8'h1F;
                    16'h021E: data_out = 8'h20;
                    16'h021F: data_out = 8'h21;
                    16'h0220: data_out = 8'h22;
                    16'h0221: data_out = 8'h23;
                    16'h0222: data_out = 8'h24;
                    16'h0223: data_out = 8'h25;
                    16'h0224: data_out = 8'h26;
                    16'h0225: data_out = 8'h27;
                    16'h0226: data_out = 8'h28;
                    16'h0227: data_out = 8'h29;
                    16'h0228: data_out = 8'h2A;
                    16'h0229: data_out = 8'h2B;
                    16'h022A: data_out = 8'h2C;
                    16'h022B: data_out = 8'h2D;
                    16'h022C: data_out = 8'h2E;
                    16'h022D: data_out = 8'h2F;
                    16'h022E: data_out = 8'h30;
                    16'h022F: data_out = 8'h31;
                    16'h0230: data_out = 8'h32;
                    16'h0231: data_out = 8'h33;
                    16'h0232: data_out = 8'h34;
                    16'h0233: data_out = 8'h35;
                    16'h0234: data_out = 8'h36;
                    16'h0235: data_out = 8'h37;
                    16'h0236: data_out = 8'h38;
                    16'h0237: data_out = 8'h39;
                    16'h0238: data_out = 8'h3A;
                    16'h0239: data_out = 8'h3B;
                    16'h023A: data_out = 8'h3C;
                    16'h023B: data_out = 8'h3D;
                    16'h023C: data_out = 8'h3E;
                    16'h023D: data_out = 8'h3F;
                    16'h023E: data_out = 8'h40;
                    16'h023F: data_out = 8'h41;
                    16'h0240: data_out = 8'h42;
                    16'h0241: data_out = 8'h43;
                    16'h0242: data_out = 8'h44;
                    16'h0243: data_out = 8'h45;
                    16'h0244: data_out = 8'h46;
                    16'h0245: data_out = 8'h47;
                    16'h0246: data_out = 8'h48;
                    16'h0247: data_out = 8'h49;
                    16'h0248: data_out = 8'h4A;
                    16'h0249: data_out = 8'h4B;
                    16'h024A: data_out = 8'h4C;
                    16'h024B: data_out = 8'h4D;
                    16'h024C: data_out = 8'h4E;
                    16'h024D: data_out = 8'h4F;
                    16'h024E: data_out = 8'h50;
                    16'h024F: data_out = 8'h51;
                    16'h0250: data_out = 8'h52;
                    16'h0251: data_out = 8'h53;
                    16'h0252: data_out = 8'h54;
                    16'h0253: data_out = 8'h55;
                    16'h0254: data_out = 8'h56;
                    16'h0255: data_out = 8'h57;
                    16'h0256: data_out = 8'h58;
                    16'h0257: data_out = 8'h59;
                    16'h0258: data_out = 8'h5A;
                    16'h0259: data_out = 8'h5B;
                    16'h025A: data_out = 8'h5C;
                    16'h025B: data_out = 8'h5D;
                    16'h025C: data_out = 8'h5E;
                    16'h025D: data_out = 8'h5F;
                    16'h025E: data_out = 8'h60;
                    16'h025F: data_out = 8'h61;
                    16'h0260: data_out = 8'h62;
                    16'h0261: data_out = 8'h63;
                    16'h0262: data_out = 8'h64;
                    16'h0263: data_out = 8'h65;
                    16'h0264: data_out = 8'h66;
                    16'h0265: data_out = 8'h67;
                    16'h0266: data_out = 8'h68;
                    16'h0267: data_out = 8'h69;
                    16'h0268: data_out = 8'h6A;
                    16'h0269: data_out = 8'h6B;
                    16'h026A: data_out = 8'h6C;
                    16'h026B: data_out = 8'h6D;
                    16'h026C: data_out = 8'h6E;
                    16'h026D: data_out = 8'h6F;
                    16'h026E: data_out = 8'h70;
                    16'h026F: data_out = 8'h71;
                    16'h0270: data_out = 8'h72;
                    16'h0271: data_out = 8'h73;
                    16'h0272: data_out = 8'h74;
                    16'h0273: data_out = 8'h75;
                    16'h0274: data_out = 8'h76;
                    16'h0275: data_out = 8'h77;
                    16'h0276: data_out = 8'h78;
                    16'h0277: data_out = 8'h79;
                    16'h0278: data_out = 8'h7A;
                    16'h0279: data_out = 8'h7B;
                    16'h027A: data_out = 8'h7C;
                    16'h027B: data_out = 8'h7D;
                    16'h027C: data_out = 8'h7E;
                    16'h027D: data_out = 8'h7F;
                    16'h027E: data_out = 8'h80;
                    16'h027F: data_out = 8'h81;
                    16'h0280: data_out = 8'h2;
                    16'h0281: data_out = 8'h1;
                    16'h0282: data_out = 8'h0;
                    16'h0283: data_out = 8'h81;
                    16'h0284: data_out = 8'h82;
                    16'h0285: data_out = 8'h83;
                    16'h0286: data_out = 8'h84;
                    16'h0287: data_out = 8'h85;
                    16'h0288: data_out = 8'h86;
                    16'h0289: data_out = 8'h87;
                    16'h028A: data_out = 8'h88;
                    16'h028B: data_out = 8'h89;
                    16'h028C: data_out = 8'h8A;
                    16'h028D: data_out = 8'h8B;
                    16'h028E: data_out = 8'h8C;
                    16'h028F: data_out = 8'h8D;
                    16'h0290: data_out = 8'h8E;
                    16'h0291: data_out = 8'h8F;
                    16'h0292: data_out = 8'h90;
                    16'h0293: data_out = 8'h91;
                    16'h0294: data_out = 8'h92;
                    16'h0295: data_out = 8'h93;
                    16'h0296: data_out = 8'h94;
                    16'h0297: data_out = 8'h95;
                    16'h0298: data_out = 8'h96;
                    16'h0299: data_out = 8'h97;
                    16'h029A: data_out = 8'h98;
                    16'h029B: data_out = 8'h99;
                    16'h029C: data_out = 8'h9A;
                    16'h029D: data_out = 8'h9B;
                    16'h029E: data_out = 8'h9C;
                    16'h029F: data_out = 8'h9D;
                    16'h02A0: data_out = 8'h9E;
                    16'h02A1: data_out = 8'h9F;
                    16'h02A2: data_out = 8'hA0;
                    16'h02A3: data_out = 8'hA1;
                    16'h02A4: data_out = 8'hA2;
                    16'h02A5: data_out = 8'hA3;
                    16'h02A6: data_out = 8'hA4;
                    16'h02A7: data_out = 8'hA5;
                    16'h02A8: data_out = 8'hA6;
                    16'h02A9: data_out = 8'hA7;
                    16'h02AA: data_out = 8'hA8;
                    16'h02AB: data_out = 8'hA9;
                    16'h02AC: data_out = 8'hAA;
                    16'h02AD: data_out = 8'hAB;
                    16'h02AE: data_out = 8'hAC;
                    16'h02AF: data_out = 8'hAD;
                    16'h02B0: data_out = 8'hAE;
                    16'h02B1: data_out = 8'hAF;
                    16'h02B2: data_out = 8'hB0;
                    16'h02B3: data_out = 8'hB1;
                    16'h02B4: data_out = 8'hB2;
                    16'h02B5: data_out = 8'hB3;
                    16'h02B6: data_out = 8'hB4;
                    16'h02B7: data_out = 8'hB5;
                    16'h02B8: data_out = 8'hB6;
                    16'h02B9: data_out = 8'hB7;
                    16'h02BA: data_out = 8'hB8;
                    16'h02BB: data_out = 8'hB9;
                    16'h02BC: data_out = 8'hBA;
                    16'h02BD: data_out = 8'hBB;
                    16'h02BE: data_out = 8'hBC;
                    16'h02BF: data_out = 8'hBD;
                    16'h02C0: data_out = 8'hBE;
                    16'h02C1: data_out = 8'hBF;
                    16'h02C2: data_out = 8'hC0;
                    16'h02C3: data_out = 8'hC1;
                    16'h02C4: data_out = 8'hC2;
                    16'h02C5: data_out = 8'hC3;
                    16'h02C6: data_out = 8'hC4;
                    16'h02C7: data_out = 8'hC5;
                    16'h02C8: data_out = 8'hC6;
                    16'h02C9: data_out = 8'hC7;
                    16'h02CA: data_out = 8'hC8;
                    16'h02CB: data_out = 8'hC9;
                    16'h02CC: data_out = 8'hCA;
                    16'h02CD: data_out = 8'hCB;
                    16'h02CE: data_out = 8'hCC;
                    16'h02CF: data_out = 8'hCD;
                    16'h02D0: data_out = 8'hCE;
                    16'h02D1: data_out = 8'hCF;
                    16'h02D2: data_out = 8'hD0;
                    16'h02D3: data_out = 8'hD1;
                    16'h02D4: data_out = 8'hD2;
                    16'h02D5: data_out = 8'hD3;
                    16'h02D6: data_out = 8'hD4;
                    16'h02D7: data_out = 8'hD5;
                    16'h02D8: data_out = 8'hD6;
                    16'h02D9: data_out = 8'hD7;
                    16'h02DA: data_out = 8'hD8;
                    16'h02DB: data_out = 8'hD9;
                    16'h02DC: data_out = 8'hDA;
                    16'h02DD: data_out = 8'hDB;
                    16'h02DE: data_out = 8'hDC;
                    16'h02DF: data_out = 8'hDD;
                    16'h02E0: data_out = 8'hDE;
                    16'h02E1: data_out = 8'hDF;
                    16'h02E2: data_out = 8'hE0;
                    16'h02E3: data_out = 8'hE1;
                    16'h02E4: data_out = 8'hE2;
                    16'h02E5: data_out = 8'hE3;
                    16'h02E6: data_out = 8'hE4;
                    16'h02E7: data_out = 8'hE5;
                    16'h02E8: data_out = 8'hE6;
                    16'h02E9: data_out = 8'hE7;
                    16'h02EA: data_out = 8'hE8;
                    16'h02EB: data_out = 8'hE9;
                    16'h02EC: data_out = 8'hEA;
                    16'h02ED: data_out = 8'hEB;
                    16'h02EE: data_out = 8'hEC;
                    16'h02EF: data_out = 8'hED;
                    16'h02F0: data_out = 8'hEE;
                    16'h02F1: data_out = 8'hEF;
                    16'h02F2: data_out = 8'hF0;
                    16'h02F3: data_out = 8'hF1;
                    16'h02F4: data_out = 8'hF2;
                    16'h02F5: data_out = 8'hF3;
                    16'h02F6: data_out = 8'hF4;
                    16'h02F7: data_out = 8'hF5;
                    16'h02F8: data_out = 8'hF6;
                    16'h02F9: data_out = 8'hF7;
                    16'h02FA: data_out = 8'hF8;
                    16'h02FB: data_out = 8'hF9;
                    16'h02FC: data_out = 8'hFA;
                    16'h02FD: data_out = 8'hFB;
                    16'h02FE: data_out = 8'hFC;
                    16'h02FF: data_out = 8'hFD;
                    16'h0300: data_out = 8'h3;
                    16'h0301: data_out = 8'h4;
                    16'h0302: data_out = 8'h5;
                    16'h0303: data_out = 8'h6;
                    16'h0304: data_out = 8'h7;
                    16'h0305: data_out = 8'h8;
                    16'h0306: data_out = 8'h9;
                    16'h0307: data_out = 8'hA;
                    16'h0308: data_out = 8'hB;
                    16'h0309: data_out = 8'hC;
                    16'h030A: data_out = 8'hD;
                    16'h030B: data_out = 8'hE;
                    16'h030C: data_out = 8'hF;
                    16'h030D: data_out = 8'h10;
                    16'h030E: data_out = 8'h11;
                    16'h030F: data_out = 8'h12;
                    16'h0310: data_out = 8'h13;
                    16'h0311: data_out = 8'h14;
                    16'h0312: data_out = 8'h15;
                    16'h0313: data_out = 8'h16;
                    16'h0314: data_out = 8'h17;
                    16'h0315: data_out = 8'h18;
                    16'h0316: data_out = 8'h19;
                    16'h0317: data_out = 8'h1A;
                    16'h0318: data_out = 8'h1B;
                    16'h0319: data_out = 8'h1C;
                    16'h031A: data_out = 8'h1D;
                    16'h031B: data_out = 8'h1E;
                    16'h031C: data_out = 8'h1F;
                    16'h031D: data_out = 8'h20;
                    16'h031E: data_out = 8'h21;
                    16'h031F: data_out = 8'h22;
                    16'h0320: data_out = 8'h23;
                    16'h0321: data_out = 8'h24;
                    16'h0322: data_out = 8'h25;
                    16'h0323: data_out = 8'h26;
                    16'h0324: data_out = 8'h27;
                    16'h0325: data_out = 8'h28;
                    16'h0326: data_out = 8'h29;
                    16'h0327: data_out = 8'h2A;
                    16'h0328: data_out = 8'h2B;
                    16'h0329: data_out = 8'h2C;
                    16'h032A: data_out = 8'h2D;
                    16'h032B: data_out = 8'h2E;
                    16'h032C: data_out = 8'h2F;
                    16'h032D: data_out = 8'h30;
                    16'h032E: data_out = 8'h31;
                    16'h032F: data_out = 8'h32;
                    16'h0330: data_out = 8'h33;
                    16'h0331: data_out = 8'h34;
                    16'h0332: data_out = 8'h35;
                    16'h0333: data_out = 8'h36;
                    16'h0334: data_out = 8'h37;
                    16'h0335: data_out = 8'h38;
                    16'h0336: data_out = 8'h39;
                    16'h0337: data_out = 8'h3A;
                    16'h0338: data_out = 8'h3B;
                    16'h0339: data_out = 8'h3C;
                    16'h033A: data_out = 8'h3D;
                    16'h033B: data_out = 8'h3E;
                    16'h033C: data_out = 8'h3F;
                    16'h033D: data_out = 8'h40;
                    16'h033E: data_out = 8'h41;
                    16'h033F: data_out = 8'h42;
                    16'h0340: data_out = 8'h43;
                    16'h0341: data_out = 8'h44;
                    16'h0342: data_out = 8'h45;
                    16'h0343: data_out = 8'h46;
                    16'h0344: data_out = 8'h47;
                    16'h0345: data_out = 8'h48;
                    16'h0346: data_out = 8'h49;
                    16'h0347: data_out = 8'h4A;
                    16'h0348: data_out = 8'h4B;
                    16'h0349: data_out = 8'h4C;
                    16'h034A: data_out = 8'h4D;
                    16'h034B: data_out = 8'h4E;
                    16'h034C: data_out = 8'h4F;
                    16'h034D: data_out = 8'h50;
                    16'h034E: data_out = 8'h51;
                    16'h034F: data_out = 8'h52;
                    16'h0350: data_out = 8'h53;
                    16'h0351: data_out = 8'h54;
                    16'h0352: data_out = 8'h55;
                    16'h0353: data_out = 8'h56;
                    16'h0354: data_out = 8'h57;
                    16'h0355: data_out = 8'h58;
                    16'h0356: data_out = 8'h59;
                    16'h0357: data_out = 8'h5A;
                    16'h0358: data_out = 8'h5B;
                    16'h0359: data_out = 8'h5C;
                    16'h035A: data_out = 8'h5D;
                    16'h035B: data_out = 8'h5E;
                    16'h035C: data_out = 8'h5F;
                    16'h035D: data_out = 8'h60;
                    16'h035E: data_out = 8'h61;
                    16'h035F: data_out = 8'h62;
                    16'h0360: data_out = 8'h63;
                    16'h0361: data_out = 8'h64;
                    16'h0362: data_out = 8'h65;
                    16'h0363: data_out = 8'h66;
                    16'h0364: data_out = 8'h67;
                    16'h0365: data_out = 8'h68;
                    16'h0366: data_out = 8'h69;
                    16'h0367: data_out = 8'h6A;
                    16'h0368: data_out = 8'h6B;
                    16'h0369: data_out = 8'h6C;
                    16'h036A: data_out = 8'h6D;
                    16'h036B: data_out = 8'h6E;
                    16'h036C: data_out = 8'h6F;
                    16'h036D: data_out = 8'h70;
                    16'h036E: data_out = 8'h71;
                    16'h036F: data_out = 8'h72;
                    16'h0370: data_out = 8'h73;
                    16'h0371: data_out = 8'h74;
                    16'h0372: data_out = 8'h75;
                    16'h0373: data_out = 8'h76;
                    16'h0374: data_out = 8'h77;
                    16'h0375: data_out = 8'h78;
                    16'h0376: data_out = 8'h79;
                    16'h0377: data_out = 8'h7A;
                    16'h0378: data_out = 8'h7B;
                    16'h0379: data_out = 8'h7C;
                    16'h037A: data_out = 8'h7D;
                    16'h037B: data_out = 8'h7E;
                    16'h037C: data_out = 8'h7F;
                    16'h037D: data_out = 8'h80;
                    16'h037E: data_out = 8'h81;
                    16'h037F: data_out = 8'h82;
                    16'h0380: data_out = 8'h3;
                    16'h0381: data_out = 8'h2;
                    16'h0382: data_out = 8'h1;
                    16'h0383: data_out = 8'h0;
                    16'h0384: data_out = 8'h81;
                    16'h0385: data_out = 8'h82;
                    16'h0386: data_out = 8'h83;
                    16'h0387: data_out = 8'h84;
                    16'h0388: data_out = 8'h85;
                    16'h0389: data_out = 8'h86;
                    16'h038A: data_out = 8'h87;
                    16'h038B: data_out = 8'h88;
                    16'h038C: data_out = 8'h89;
                    16'h038D: data_out = 8'h8A;
                    16'h038E: data_out = 8'h8B;
                    16'h038F: data_out = 8'h8C;
                    16'h0390: data_out = 8'h8D;
                    16'h0391: data_out = 8'h8E;
                    16'h0392: data_out = 8'h8F;
                    16'h0393: data_out = 8'h90;
                    16'h0394: data_out = 8'h91;
                    16'h0395: data_out = 8'h92;
                    16'h0396: data_out = 8'h93;
                    16'h0397: data_out = 8'h94;
                    16'h0398: data_out = 8'h95;
                    16'h0399: data_out = 8'h96;
                    16'h039A: data_out = 8'h97;
                    16'h039B: data_out = 8'h98;
                    16'h039C: data_out = 8'h99;
                    16'h039D: data_out = 8'h9A;
                    16'h039E: data_out = 8'h9B;
                    16'h039F: data_out = 8'h9C;
                    16'h03A0: data_out = 8'h9D;
                    16'h03A1: data_out = 8'h9E;
                    16'h03A2: data_out = 8'h9F;
                    16'h03A3: data_out = 8'hA0;
                    16'h03A4: data_out = 8'hA1;
                    16'h03A5: data_out = 8'hA2;
                    16'h03A6: data_out = 8'hA3;
                    16'h03A7: data_out = 8'hA4;
                    16'h03A8: data_out = 8'hA5;
                    16'h03A9: data_out = 8'hA6;
                    16'h03AA: data_out = 8'hA7;
                    16'h03AB: data_out = 8'hA8;
                    16'h03AC: data_out = 8'hA9;
                    16'h03AD: data_out = 8'hAA;
                    16'h03AE: data_out = 8'hAB;
                    16'h03AF: data_out = 8'hAC;
                    16'h03B0: data_out = 8'hAD;
                    16'h03B1: data_out = 8'hAE;
                    16'h03B2: data_out = 8'hAF;
                    16'h03B3: data_out = 8'hB0;
                    16'h03B4: data_out = 8'hB1;
                    16'h03B5: data_out = 8'hB2;
                    16'h03B6: data_out = 8'hB3;
                    16'h03B7: data_out = 8'hB4;
                    16'h03B8: data_out = 8'hB5;
                    16'h03B9: data_out = 8'hB6;
                    16'h03BA: data_out = 8'hB7;
                    16'h03BB: data_out = 8'hB8;
                    16'h03BC: data_out = 8'hB9;
                    16'h03BD: data_out = 8'hBA;
                    16'h03BE: data_out = 8'hBB;
                    16'h03BF: data_out = 8'hBC;
                    16'h03C0: data_out = 8'hBD;
                    16'h03C1: data_out = 8'hBE;
                    16'h03C2: data_out = 8'hBF;
                    16'h03C3: data_out = 8'hC0;
                    16'h03C4: data_out = 8'hC1;
                    16'h03C5: data_out = 8'hC2;
                    16'h03C6: data_out = 8'hC3;
                    16'h03C7: data_out = 8'hC4;
                    16'h03C8: data_out = 8'hC5;
                    16'h03C9: data_out = 8'hC6;
                    16'h03CA: data_out = 8'hC7;
                    16'h03CB: data_out = 8'hC8;
                    16'h03CC: data_out = 8'hC9;
                    16'h03CD: data_out = 8'hCA;
                    16'h03CE: data_out = 8'hCB;
                    16'h03CF: data_out = 8'hCC;
                    16'h03D0: data_out = 8'hCD;
                    16'h03D1: data_out = 8'hCE;
                    16'h03D2: data_out = 8'hCF;
                    16'h03D3: data_out = 8'hD0;
                    16'h03D4: data_out = 8'hD1;
                    16'h03D5: data_out = 8'hD2;
                    16'h03D6: data_out = 8'hD3;
                    16'h03D7: data_out = 8'hD4;
                    16'h03D8: data_out = 8'hD5;
                    16'h03D9: data_out = 8'hD6;
                    16'h03DA: data_out = 8'hD7;
                    16'h03DB: data_out = 8'hD8;
                    16'h03DC: data_out = 8'hD9;
                    16'h03DD: data_out = 8'hDA;
                    16'h03DE: data_out = 8'hDB;
                    16'h03DF: data_out = 8'hDC;
                    16'h03E0: data_out = 8'hDD;
                    16'h03E1: data_out = 8'hDE;
                    16'h03E2: data_out = 8'hDF;
                    16'h03E3: data_out = 8'hE0;
                    16'h03E4: data_out = 8'hE1;
                    16'h03E5: data_out = 8'hE2;
                    16'h03E6: data_out = 8'hE3;
                    16'h03E7: data_out = 8'hE4;
                    16'h03E8: data_out = 8'hE5;
                    16'h03E9: data_out = 8'hE6;
                    16'h03EA: data_out = 8'hE7;
                    16'h03EB: data_out = 8'hE8;
                    16'h03EC: data_out = 8'hE9;
                    16'h03ED: data_out = 8'hEA;
                    16'h03EE: data_out = 8'hEB;
                    16'h03EF: data_out = 8'hEC;
                    16'h03F0: data_out = 8'hED;
                    16'h03F1: data_out = 8'hEE;
                    16'h03F2: data_out = 8'hEF;
                    16'h03F3: data_out = 8'hF0;
                    16'h03F4: data_out = 8'hF1;
                    16'h03F5: data_out = 8'hF2;
                    16'h03F6: data_out = 8'hF3;
                    16'h03F7: data_out = 8'hF4;
                    16'h03F8: data_out = 8'hF5;
                    16'h03F9: data_out = 8'hF6;
                    16'h03FA: data_out = 8'hF7;
                    16'h03FB: data_out = 8'hF8;
                    16'h03FC: data_out = 8'hF9;
                    16'h03FD: data_out = 8'hFA;
                    16'h03FE: data_out = 8'hFB;
                    16'h03FF: data_out = 8'hFC;
                    16'h0400: data_out = 8'h4;
                    16'h0401: data_out = 8'h5;
                    16'h0402: data_out = 8'h6;
                    16'h0403: data_out = 8'h7;
                    16'h0404: data_out = 8'h8;
                    16'h0405: data_out = 8'h9;
                    16'h0406: data_out = 8'hA;
                    16'h0407: data_out = 8'hB;
                    16'h0408: data_out = 8'hC;
                    16'h0409: data_out = 8'hD;
                    16'h040A: data_out = 8'hE;
                    16'h040B: data_out = 8'hF;
                    16'h040C: data_out = 8'h10;
                    16'h040D: data_out = 8'h11;
                    16'h040E: data_out = 8'h12;
                    16'h040F: data_out = 8'h13;
                    16'h0410: data_out = 8'h14;
                    16'h0411: data_out = 8'h15;
                    16'h0412: data_out = 8'h16;
                    16'h0413: data_out = 8'h17;
                    16'h0414: data_out = 8'h18;
                    16'h0415: data_out = 8'h19;
                    16'h0416: data_out = 8'h1A;
                    16'h0417: data_out = 8'h1B;
                    16'h0418: data_out = 8'h1C;
                    16'h0419: data_out = 8'h1D;
                    16'h041A: data_out = 8'h1E;
                    16'h041B: data_out = 8'h1F;
                    16'h041C: data_out = 8'h20;
                    16'h041D: data_out = 8'h21;
                    16'h041E: data_out = 8'h22;
                    16'h041F: data_out = 8'h23;
                    16'h0420: data_out = 8'h24;
                    16'h0421: data_out = 8'h25;
                    16'h0422: data_out = 8'h26;
                    16'h0423: data_out = 8'h27;
                    16'h0424: data_out = 8'h28;
                    16'h0425: data_out = 8'h29;
                    16'h0426: data_out = 8'h2A;
                    16'h0427: data_out = 8'h2B;
                    16'h0428: data_out = 8'h2C;
                    16'h0429: data_out = 8'h2D;
                    16'h042A: data_out = 8'h2E;
                    16'h042B: data_out = 8'h2F;
                    16'h042C: data_out = 8'h30;
                    16'h042D: data_out = 8'h31;
                    16'h042E: data_out = 8'h32;
                    16'h042F: data_out = 8'h33;
                    16'h0430: data_out = 8'h34;
                    16'h0431: data_out = 8'h35;
                    16'h0432: data_out = 8'h36;
                    16'h0433: data_out = 8'h37;
                    16'h0434: data_out = 8'h38;
                    16'h0435: data_out = 8'h39;
                    16'h0436: data_out = 8'h3A;
                    16'h0437: data_out = 8'h3B;
                    16'h0438: data_out = 8'h3C;
                    16'h0439: data_out = 8'h3D;
                    16'h043A: data_out = 8'h3E;
                    16'h043B: data_out = 8'h3F;
                    16'h043C: data_out = 8'h40;
                    16'h043D: data_out = 8'h41;
                    16'h043E: data_out = 8'h42;
                    16'h043F: data_out = 8'h43;
                    16'h0440: data_out = 8'h44;
                    16'h0441: data_out = 8'h45;
                    16'h0442: data_out = 8'h46;
                    16'h0443: data_out = 8'h47;
                    16'h0444: data_out = 8'h48;
                    16'h0445: data_out = 8'h49;
                    16'h0446: data_out = 8'h4A;
                    16'h0447: data_out = 8'h4B;
                    16'h0448: data_out = 8'h4C;
                    16'h0449: data_out = 8'h4D;
                    16'h044A: data_out = 8'h4E;
                    16'h044B: data_out = 8'h4F;
                    16'h044C: data_out = 8'h50;
                    16'h044D: data_out = 8'h51;
                    16'h044E: data_out = 8'h52;
                    16'h044F: data_out = 8'h53;
                    16'h0450: data_out = 8'h54;
                    16'h0451: data_out = 8'h55;
                    16'h0452: data_out = 8'h56;
                    16'h0453: data_out = 8'h57;
                    16'h0454: data_out = 8'h58;
                    16'h0455: data_out = 8'h59;
                    16'h0456: data_out = 8'h5A;
                    16'h0457: data_out = 8'h5B;
                    16'h0458: data_out = 8'h5C;
                    16'h0459: data_out = 8'h5D;
                    16'h045A: data_out = 8'h5E;
                    16'h045B: data_out = 8'h5F;
                    16'h045C: data_out = 8'h60;
                    16'h045D: data_out = 8'h61;
                    16'h045E: data_out = 8'h62;
                    16'h045F: data_out = 8'h63;
                    16'h0460: data_out = 8'h64;
                    16'h0461: data_out = 8'h65;
                    16'h0462: data_out = 8'h66;
                    16'h0463: data_out = 8'h67;
                    16'h0464: data_out = 8'h68;
                    16'h0465: data_out = 8'h69;
                    16'h0466: data_out = 8'h6A;
                    16'h0467: data_out = 8'h6B;
                    16'h0468: data_out = 8'h6C;
                    16'h0469: data_out = 8'h6D;
                    16'h046A: data_out = 8'h6E;
                    16'h046B: data_out = 8'h6F;
                    16'h046C: data_out = 8'h70;
                    16'h046D: data_out = 8'h71;
                    16'h046E: data_out = 8'h72;
                    16'h046F: data_out = 8'h73;
                    16'h0470: data_out = 8'h74;
                    16'h0471: data_out = 8'h75;
                    16'h0472: data_out = 8'h76;
                    16'h0473: data_out = 8'h77;
                    16'h0474: data_out = 8'h78;
                    16'h0475: data_out = 8'h79;
                    16'h0476: data_out = 8'h7A;
                    16'h0477: data_out = 8'h7B;
                    16'h0478: data_out = 8'h7C;
                    16'h0479: data_out = 8'h7D;
                    16'h047A: data_out = 8'h7E;
                    16'h047B: data_out = 8'h7F;
                    16'h047C: data_out = 8'h80;
                    16'h047D: data_out = 8'h81;
                    16'h047E: data_out = 8'h82;
                    16'h047F: data_out = 8'h83;
                    16'h0480: data_out = 8'h4;
                    16'h0481: data_out = 8'h3;
                    16'h0482: data_out = 8'h2;
                    16'h0483: data_out = 8'h1;
                    16'h0484: data_out = 8'h0;
                    16'h0485: data_out = 8'h81;
                    16'h0486: data_out = 8'h82;
                    16'h0487: data_out = 8'h83;
                    16'h0488: data_out = 8'h84;
                    16'h0489: data_out = 8'h85;
                    16'h048A: data_out = 8'h86;
                    16'h048B: data_out = 8'h87;
                    16'h048C: data_out = 8'h88;
                    16'h048D: data_out = 8'h89;
                    16'h048E: data_out = 8'h8A;
                    16'h048F: data_out = 8'h8B;
                    16'h0490: data_out = 8'h8C;
                    16'h0491: data_out = 8'h8D;
                    16'h0492: data_out = 8'h8E;
                    16'h0493: data_out = 8'h8F;
                    16'h0494: data_out = 8'h90;
                    16'h0495: data_out = 8'h91;
                    16'h0496: data_out = 8'h92;
                    16'h0497: data_out = 8'h93;
                    16'h0498: data_out = 8'h94;
                    16'h0499: data_out = 8'h95;
                    16'h049A: data_out = 8'h96;
                    16'h049B: data_out = 8'h97;
                    16'h049C: data_out = 8'h98;
                    16'h049D: data_out = 8'h99;
                    16'h049E: data_out = 8'h9A;
                    16'h049F: data_out = 8'h9B;
                    16'h04A0: data_out = 8'h9C;
                    16'h04A1: data_out = 8'h9D;
                    16'h04A2: data_out = 8'h9E;
                    16'h04A3: data_out = 8'h9F;
                    16'h04A4: data_out = 8'hA0;
                    16'h04A5: data_out = 8'hA1;
                    16'h04A6: data_out = 8'hA2;
                    16'h04A7: data_out = 8'hA3;
                    16'h04A8: data_out = 8'hA4;
                    16'h04A9: data_out = 8'hA5;
                    16'h04AA: data_out = 8'hA6;
                    16'h04AB: data_out = 8'hA7;
                    16'h04AC: data_out = 8'hA8;
                    16'h04AD: data_out = 8'hA9;
                    16'h04AE: data_out = 8'hAA;
                    16'h04AF: data_out = 8'hAB;
                    16'h04B0: data_out = 8'hAC;
                    16'h04B1: data_out = 8'hAD;
                    16'h04B2: data_out = 8'hAE;
                    16'h04B3: data_out = 8'hAF;
                    16'h04B4: data_out = 8'hB0;
                    16'h04B5: data_out = 8'hB1;
                    16'h04B6: data_out = 8'hB2;
                    16'h04B7: data_out = 8'hB3;
                    16'h04B8: data_out = 8'hB4;
                    16'h04B9: data_out = 8'hB5;
                    16'h04BA: data_out = 8'hB6;
                    16'h04BB: data_out = 8'hB7;
                    16'h04BC: data_out = 8'hB8;
                    16'h04BD: data_out = 8'hB9;
                    16'h04BE: data_out = 8'hBA;
                    16'h04BF: data_out = 8'hBB;
                    16'h04C0: data_out = 8'hBC;
                    16'h04C1: data_out = 8'hBD;
                    16'h04C2: data_out = 8'hBE;
                    16'h04C3: data_out = 8'hBF;
                    16'h04C4: data_out = 8'hC0;
                    16'h04C5: data_out = 8'hC1;
                    16'h04C6: data_out = 8'hC2;
                    16'h04C7: data_out = 8'hC3;
                    16'h04C8: data_out = 8'hC4;
                    16'h04C9: data_out = 8'hC5;
                    16'h04CA: data_out = 8'hC6;
                    16'h04CB: data_out = 8'hC7;
                    16'h04CC: data_out = 8'hC8;
                    16'h04CD: data_out = 8'hC9;
                    16'h04CE: data_out = 8'hCA;
                    16'h04CF: data_out = 8'hCB;
                    16'h04D0: data_out = 8'hCC;
                    16'h04D1: data_out = 8'hCD;
                    16'h04D2: data_out = 8'hCE;
                    16'h04D3: data_out = 8'hCF;
                    16'h04D4: data_out = 8'hD0;
                    16'h04D5: data_out = 8'hD1;
                    16'h04D6: data_out = 8'hD2;
                    16'h04D7: data_out = 8'hD3;
                    16'h04D8: data_out = 8'hD4;
                    16'h04D9: data_out = 8'hD5;
                    16'h04DA: data_out = 8'hD6;
                    16'h04DB: data_out = 8'hD7;
                    16'h04DC: data_out = 8'hD8;
                    16'h04DD: data_out = 8'hD9;
                    16'h04DE: data_out = 8'hDA;
                    16'h04DF: data_out = 8'hDB;
                    16'h04E0: data_out = 8'hDC;
                    16'h04E1: data_out = 8'hDD;
                    16'h04E2: data_out = 8'hDE;
                    16'h04E3: data_out = 8'hDF;
                    16'h04E4: data_out = 8'hE0;
                    16'h04E5: data_out = 8'hE1;
                    16'h04E6: data_out = 8'hE2;
                    16'h04E7: data_out = 8'hE3;
                    16'h04E8: data_out = 8'hE4;
                    16'h04E9: data_out = 8'hE5;
                    16'h04EA: data_out = 8'hE6;
                    16'h04EB: data_out = 8'hE7;
                    16'h04EC: data_out = 8'hE8;
                    16'h04ED: data_out = 8'hE9;
                    16'h04EE: data_out = 8'hEA;
                    16'h04EF: data_out = 8'hEB;
                    16'h04F0: data_out = 8'hEC;
                    16'h04F1: data_out = 8'hED;
                    16'h04F2: data_out = 8'hEE;
                    16'h04F3: data_out = 8'hEF;
                    16'h04F4: data_out = 8'hF0;
                    16'h04F5: data_out = 8'hF1;
                    16'h04F6: data_out = 8'hF2;
                    16'h04F7: data_out = 8'hF3;
                    16'h04F8: data_out = 8'hF4;
                    16'h04F9: data_out = 8'hF5;
                    16'h04FA: data_out = 8'hF6;
                    16'h04FB: data_out = 8'hF7;
                    16'h04FC: data_out = 8'hF8;
                    16'h04FD: data_out = 8'hF9;
                    16'h04FE: data_out = 8'hFA;
                    16'h04FF: data_out = 8'hFB;
                    16'h0500: data_out = 8'h5;
                    16'h0501: data_out = 8'h6;
                    16'h0502: data_out = 8'h7;
                    16'h0503: data_out = 8'h8;
                    16'h0504: data_out = 8'h9;
                    16'h0505: data_out = 8'hA;
                    16'h0506: data_out = 8'hB;
                    16'h0507: data_out = 8'hC;
                    16'h0508: data_out = 8'hD;
                    16'h0509: data_out = 8'hE;
                    16'h050A: data_out = 8'hF;
                    16'h050B: data_out = 8'h10;
                    16'h050C: data_out = 8'h11;
                    16'h050D: data_out = 8'h12;
                    16'h050E: data_out = 8'h13;
                    16'h050F: data_out = 8'h14;
                    16'h0510: data_out = 8'h15;
                    16'h0511: data_out = 8'h16;
                    16'h0512: data_out = 8'h17;
                    16'h0513: data_out = 8'h18;
                    16'h0514: data_out = 8'h19;
                    16'h0515: data_out = 8'h1A;
                    16'h0516: data_out = 8'h1B;
                    16'h0517: data_out = 8'h1C;
                    16'h0518: data_out = 8'h1D;
                    16'h0519: data_out = 8'h1E;
                    16'h051A: data_out = 8'h1F;
                    16'h051B: data_out = 8'h20;
                    16'h051C: data_out = 8'h21;
                    16'h051D: data_out = 8'h22;
                    16'h051E: data_out = 8'h23;
                    16'h051F: data_out = 8'h24;
                    16'h0520: data_out = 8'h25;
                    16'h0521: data_out = 8'h26;
                    16'h0522: data_out = 8'h27;
                    16'h0523: data_out = 8'h28;
                    16'h0524: data_out = 8'h29;
                    16'h0525: data_out = 8'h2A;
                    16'h0526: data_out = 8'h2B;
                    16'h0527: data_out = 8'h2C;
                    16'h0528: data_out = 8'h2D;
                    16'h0529: data_out = 8'h2E;
                    16'h052A: data_out = 8'h2F;
                    16'h052B: data_out = 8'h30;
                    16'h052C: data_out = 8'h31;
                    16'h052D: data_out = 8'h32;
                    16'h052E: data_out = 8'h33;
                    16'h052F: data_out = 8'h34;
                    16'h0530: data_out = 8'h35;
                    16'h0531: data_out = 8'h36;
                    16'h0532: data_out = 8'h37;
                    16'h0533: data_out = 8'h38;
                    16'h0534: data_out = 8'h39;
                    16'h0535: data_out = 8'h3A;
                    16'h0536: data_out = 8'h3B;
                    16'h0537: data_out = 8'h3C;
                    16'h0538: data_out = 8'h3D;
                    16'h0539: data_out = 8'h3E;
                    16'h053A: data_out = 8'h3F;
                    16'h053B: data_out = 8'h40;
                    16'h053C: data_out = 8'h41;
                    16'h053D: data_out = 8'h42;
                    16'h053E: data_out = 8'h43;
                    16'h053F: data_out = 8'h44;
                    16'h0540: data_out = 8'h45;
                    16'h0541: data_out = 8'h46;
                    16'h0542: data_out = 8'h47;
                    16'h0543: data_out = 8'h48;
                    16'h0544: data_out = 8'h49;
                    16'h0545: data_out = 8'h4A;
                    16'h0546: data_out = 8'h4B;
                    16'h0547: data_out = 8'h4C;
                    16'h0548: data_out = 8'h4D;
                    16'h0549: data_out = 8'h4E;
                    16'h054A: data_out = 8'h4F;
                    16'h054B: data_out = 8'h50;
                    16'h054C: data_out = 8'h51;
                    16'h054D: data_out = 8'h52;
                    16'h054E: data_out = 8'h53;
                    16'h054F: data_out = 8'h54;
                    16'h0550: data_out = 8'h55;
                    16'h0551: data_out = 8'h56;
                    16'h0552: data_out = 8'h57;
                    16'h0553: data_out = 8'h58;
                    16'h0554: data_out = 8'h59;
                    16'h0555: data_out = 8'h5A;
                    16'h0556: data_out = 8'h5B;
                    16'h0557: data_out = 8'h5C;
                    16'h0558: data_out = 8'h5D;
                    16'h0559: data_out = 8'h5E;
                    16'h055A: data_out = 8'h5F;
                    16'h055B: data_out = 8'h60;
                    16'h055C: data_out = 8'h61;
                    16'h055D: data_out = 8'h62;
                    16'h055E: data_out = 8'h63;
                    16'h055F: data_out = 8'h64;
                    16'h0560: data_out = 8'h65;
                    16'h0561: data_out = 8'h66;
                    16'h0562: data_out = 8'h67;
                    16'h0563: data_out = 8'h68;
                    16'h0564: data_out = 8'h69;
                    16'h0565: data_out = 8'h6A;
                    16'h0566: data_out = 8'h6B;
                    16'h0567: data_out = 8'h6C;
                    16'h0568: data_out = 8'h6D;
                    16'h0569: data_out = 8'h6E;
                    16'h056A: data_out = 8'h6F;
                    16'h056B: data_out = 8'h70;
                    16'h056C: data_out = 8'h71;
                    16'h056D: data_out = 8'h72;
                    16'h056E: data_out = 8'h73;
                    16'h056F: data_out = 8'h74;
                    16'h0570: data_out = 8'h75;
                    16'h0571: data_out = 8'h76;
                    16'h0572: data_out = 8'h77;
                    16'h0573: data_out = 8'h78;
                    16'h0574: data_out = 8'h79;
                    16'h0575: data_out = 8'h7A;
                    16'h0576: data_out = 8'h7B;
                    16'h0577: data_out = 8'h7C;
                    16'h0578: data_out = 8'h7D;
                    16'h0579: data_out = 8'h7E;
                    16'h057A: data_out = 8'h7F;
                    16'h057B: data_out = 8'h80;
                    16'h057C: data_out = 8'h81;
                    16'h057D: data_out = 8'h82;
                    16'h057E: data_out = 8'h83;
                    16'h057F: data_out = 8'h84;
                    16'h0580: data_out = 8'h5;
                    16'h0581: data_out = 8'h4;
                    16'h0582: data_out = 8'h3;
                    16'h0583: data_out = 8'h2;
                    16'h0584: data_out = 8'h1;
                    16'h0585: data_out = 8'h0;
                    16'h0586: data_out = 8'h81;
                    16'h0587: data_out = 8'h82;
                    16'h0588: data_out = 8'h83;
                    16'h0589: data_out = 8'h84;
                    16'h058A: data_out = 8'h85;
                    16'h058B: data_out = 8'h86;
                    16'h058C: data_out = 8'h87;
                    16'h058D: data_out = 8'h88;
                    16'h058E: data_out = 8'h89;
                    16'h058F: data_out = 8'h8A;
                    16'h0590: data_out = 8'h8B;
                    16'h0591: data_out = 8'h8C;
                    16'h0592: data_out = 8'h8D;
                    16'h0593: data_out = 8'h8E;
                    16'h0594: data_out = 8'h8F;
                    16'h0595: data_out = 8'h90;
                    16'h0596: data_out = 8'h91;
                    16'h0597: data_out = 8'h92;
                    16'h0598: data_out = 8'h93;
                    16'h0599: data_out = 8'h94;
                    16'h059A: data_out = 8'h95;
                    16'h059B: data_out = 8'h96;
                    16'h059C: data_out = 8'h97;
                    16'h059D: data_out = 8'h98;
                    16'h059E: data_out = 8'h99;
                    16'h059F: data_out = 8'h9A;
                    16'h05A0: data_out = 8'h9B;
                    16'h05A1: data_out = 8'h9C;
                    16'h05A2: data_out = 8'h9D;
                    16'h05A3: data_out = 8'h9E;
                    16'h05A4: data_out = 8'h9F;
                    16'h05A5: data_out = 8'hA0;
                    16'h05A6: data_out = 8'hA1;
                    16'h05A7: data_out = 8'hA2;
                    16'h05A8: data_out = 8'hA3;
                    16'h05A9: data_out = 8'hA4;
                    16'h05AA: data_out = 8'hA5;
                    16'h05AB: data_out = 8'hA6;
                    16'h05AC: data_out = 8'hA7;
                    16'h05AD: data_out = 8'hA8;
                    16'h05AE: data_out = 8'hA9;
                    16'h05AF: data_out = 8'hAA;
                    16'h05B0: data_out = 8'hAB;
                    16'h05B1: data_out = 8'hAC;
                    16'h05B2: data_out = 8'hAD;
                    16'h05B3: data_out = 8'hAE;
                    16'h05B4: data_out = 8'hAF;
                    16'h05B5: data_out = 8'hB0;
                    16'h05B6: data_out = 8'hB1;
                    16'h05B7: data_out = 8'hB2;
                    16'h05B8: data_out = 8'hB3;
                    16'h05B9: data_out = 8'hB4;
                    16'h05BA: data_out = 8'hB5;
                    16'h05BB: data_out = 8'hB6;
                    16'h05BC: data_out = 8'hB7;
                    16'h05BD: data_out = 8'hB8;
                    16'h05BE: data_out = 8'hB9;
                    16'h05BF: data_out = 8'hBA;
                    16'h05C0: data_out = 8'hBB;
                    16'h05C1: data_out = 8'hBC;
                    16'h05C2: data_out = 8'hBD;
                    16'h05C3: data_out = 8'hBE;
                    16'h05C4: data_out = 8'hBF;
                    16'h05C5: data_out = 8'hC0;
                    16'h05C6: data_out = 8'hC1;
                    16'h05C7: data_out = 8'hC2;
                    16'h05C8: data_out = 8'hC3;
                    16'h05C9: data_out = 8'hC4;
                    16'h05CA: data_out = 8'hC5;
                    16'h05CB: data_out = 8'hC6;
                    16'h05CC: data_out = 8'hC7;
                    16'h05CD: data_out = 8'hC8;
                    16'h05CE: data_out = 8'hC9;
                    16'h05CF: data_out = 8'hCA;
                    16'h05D0: data_out = 8'hCB;
                    16'h05D1: data_out = 8'hCC;
                    16'h05D2: data_out = 8'hCD;
                    16'h05D3: data_out = 8'hCE;
                    16'h05D4: data_out = 8'hCF;
                    16'h05D5: data_out = 8'hD0;
                    16'h05D6: data_out = 8'hD1;
                    16'h05D7: data_out = 8'hD2;
                    16'h05D8: data_out = 8'hD3;
                    16'h05D9: data_out = 8'hD4;
                    16'h05DA: data_out = 8'hD5;
                    16'h05DB: data_out = 8'hD6;
                    16'h05DC: data_out = 8'hD7;
                    16'h05DD: data_out = 8'hD8;
                    16'h05DE: data_out = 8'hD9;
                    16'h05DF: data_out = 8'hDA;
                    16'h05E0: data_out = 8'hDB;
                    16'h05E1: data_out = 8'hDC;
                    16'h05E2: data_out = 8'hDD;
                    16'h05E3: data_out = 8'hDE;
                    16'h05E4: data_out = 8'hDF;
                    16'h05E5: data_out = 8'hE0;
                    16'h05E6: data_out = 8'hE1;
                    16'h05E7: data_out = 8'hE2;
                    16'h05E8: data_out = 8'hE3;
                    16'h05E9: data_out = 8'hE4;
                    16'h05EA: data_out = 8'hE5;
                    16'h05EB: data_out = 8'hE6;
                    16'h05EC: data_out = 8'hE7;
                    16'h05ED: data_out = 8'hE8;
                    16'h05EE: data_out = 8'hE9;
                    16'h05EF: data_out = 8'hEA;
                    16'h05F0: data_out = 8'hEB;
                    16'h05F1: data_out = 8'hEC;
                    16'h05F2: data_out = 8'hED;
                    16'h05F3: data_out = 8'hEE;
                    16'h05F4: data_out = 8'hEF;
                    16'h05F5: data_out = 8'hF0;
                    16'h05F6: data_out = 8'hF1;
                    16'h05F7: data_out = 8'hF2;
                    16'h05F8: data_out = 8'hF3;
                    16'h05F9: data_out = 8'hF4;
                    16'h05FA: data_out = 8'hF5;
                    16'h05FB: data_out = 8'hF6;
                    16'h05FC: data_out = 8'hF7;
                    16'h05FD: data_out = 8'hF8;
                    16'h05FE: data_out = 8'hF9;
                    16'h05FF: data_out = 8'hFA;
                    16'h0600: data_out = 8'h6;
                    16'h0601: data_out = 8'h7;
                    16'h0602: data_out = 8'h8;
                    16'h0603: data_out = 8'h9;
                    16'h0604: data_out = 8'hA;
                    16'h0605: data_out = 8'hB;
                    16'h0606: data_out = 8'hC;
                    16'h0607: data_out = 8'hD;
                    16'h0608: data_out = 8'hE;
                    16'h0609: data_out = 8'hF;
                    16'h060A: data_out = 8'h10;
                    16'h060B: data_out = 8'h11;
                    16'h060C: data_out = 8'h12;
                    16'h060D: data_out = 8'h13;
                    16'h060E: data_out = 8'h14;
                    16'h060F: data_out = 8'h15;
                    16'h0610: data_out = 8'h16;
                    16'h0611: data_out = 8'h17;
                    16'h0612: data_out = 8'h18;
                    16'h0613: data_out = 8'h19;
                    16'h0614: data_out = 8'h1A;
                    16'h0615: data_out = 8'h1B;
                    16'h0616: data_out = 8'h1C;
                    16'h0617: data_out = 8'h1D;
                    16'h0618: data_out = 8'h1E;
                    16'h0619: data_out = 8'h1F;
                    16'h061A: data_out = 8'h20;
                    16'h061B: data_out = 8'h21;
                    16'h061C: data_out = 8'h22;
                    16'h061D: data_out = 8'h23;
                    16'h061E: data_out = 8'h24;
                    16'h061F: data_out = 8'h25;
                    16'h0620: data_out = 8'h26;
                    16'h0621: data_out = 8'h27;
                    16'h0622: data_out = 8'h28;
                    16'h0623: data_out = 8'h29;
                    16'h0624: data_out = 8'h2A;
                    16'h0625: data_out = 8'h2B;
                    16'h0626: data_out = 8'h2C;
                    16'h0627: data_out = 8'h2D;
                    16'h0628: data_out = 8'h2E;
                    16'h0629: data_out = 8'h2F;
                    16'h062A: data_out = 8'h30;
                    16'h062B: data_out = 8'h31;
                    16'h062C: data_out = 8'h32;
                    16'h062D: data_out = 8'h33;
                    16'h062E: data_out = 8'h34;
                    16'h062F: data_out = 8'h35;
                    16'h0630: data_out = 8'h36;
                    16'h0631: data_out = 8'h37;
                    16'h0632: data_out = 8'h38;
                    16'h0633: data_out = 8'h39;
                    16'h0634: data_out = 8'h3A;
                    16'h0635: data_out = 8'h3B;
                    16'h0636: data_out = 8'h3C;
                    16'h0637: data_out = 8'h3D;
                    16'h0638: data_out = 8'h3E;
                    16'h0639: data_out = 8'h3F;
                    16'h063A: data_out = 8'h40;
                    16'h063B: data_out = 8'h41;
                    16'h063C: data_out = 8'h42;
                    16'h063D: data_out = 8'h43;
                    16'h063E: data_out = 8'h44;
                    16'h063F: data_out = 8'h45;
                    16'h0640: data_out = 8'h46;
                    16'h0641: data_out = 8'h47;
                    16'h0642: data_out = 8'h48;
                    16'h0643: data_out = 8'h49;
                    16'h0644: data_out = 8'h4A;
                    16'h0645: data_out = 8'h4B;
                    16'h0646: data_out = 8'h4C;
                    16'h0647: data_out = 8'h4D;
                    16'h0648: data_out = 8'h4E;
                    16'h0649: data_out = 8'h4F;
                    16'h064A: data_out = 8'h50;
                    16'h064B: data_out = 8'h51;
                    16'h064C: data_out = 8'h52;
                    16'h064D: data_out = 8'h53;
                    16'h064E: data_out = 8'h54;
                    16'h064F: data_out = 8'h55;
                    16'h0650: data_out = 8'h56;
                    16'h0651: data_out = 8'h57;
                    16'h0652: data_out = 8'h58;
                    16'h0653: data_out = 8'h59;
                    16'h0654: data_out = 8'h5A;
                    16'h0655: data_out = 8'h5B;
                    16'h0656: data_out = 8'h5C;
                    16'h0657: data_out = 8'h5D;
                    16'h0658: data_out = 8'h5E;
                    16'h0659: data_out = 8'h5F;
                    16'h065A: data_out = 8'h60;
                    16'h065B: data_out = 8'h61;
                    16'h065C: data_out = 8'h62;
                    16'h065D: data_out = 8'h63;
                    16'h065E: data_out = 8'h64;
                    16'h065F: data_out = 8'h65;
                    16'h0660: data_out = 8'h66;
                    16'h0661: data_out = 8'h67;
                    16'h0662: data_out = 8'h68;
                    16'h0663: data_out = 8'h69;
                    16'h0664: data_out = 8'h6A;
                    16'h0665: data_out = 8'h6B;
                    16'h0666: data_out = 8'h6C;
                    16'h0667: data_out = 8'h6D;
                    16'h0668: data_out = 8'h6E;
                    16'h0669: data_out = 8'h6F;
                    16'h066A: data_out = 8'h70;
                    16'h066B: data_out = 8'h71;
                    16'h066C: data_out = 8'h72;
                    16'h066D: data_out = 8'h73;
                    16'h066E: data_out = 8'h74;
                    16'h066F: data_out = 8'h75;
                    16'h0670: data_out = 8'h76;
                    16'h0671: data_out = 8'h77;
                    16'h0672: data_out = 8'h78;
                    16'h0673: data_out = 8'h79;
                    16'h0674: data_out = 8'h7A;
                    16'h0675: data_out = 8'h7B;
                    16'h0676: data_out = 8'h7C;
                    16'h0677: data_out = 8'h7D;
                    16'h0678: data_out = 8'h7E;
                    16'h0679: data_out = 8'h7F;
                    16'h067A: data_out = 8'h80;
                    16'h067B: data_out = 8'h81;
                    16'h067C: data_out = 8'h82;
                    16'h067D: data_out = 8'h83;
                    16'h067E: data_out = 8'h84;
                    16'h067F: data_out = 8'h85;
                    16'h0680: data_out = 8'h6;
                    16'h0681: data_out = 8'h5;
                    16'h0682: data_out = 8'h4;
                    16'h0683: data_out = 8'h3;
                    16'h0684: data_out = 8'h2;
                    16'h0685: data_out = 8'h1;
                    16'h0686: data_out = 8'h0;
                    16'h0687: data_out = 8'h81;
                    16'h0688: data_out = 8'h82;
                    16'h0689: data_out = 8'h83;
                    16'h068A: data_out = 8'h84;
                    16'h068B: data_out = 8'h85;
                    16'h068C: data_out = 8'h86;
                    16'h068D: data_out = 8'h87;
                    16'h068E: data_out = 8'h88;
                    16'h068F: data_out = 8'h89;
                    16'h0690: data_out = 8'h8A;
                    16'h0691: data_out = 8'h8B;
                    16'h0692: data_out = 8'h8C;
                    16'h0693: data_out = 8'h8D;
                    16'h0694: data_out = 8'h8E;
                    16'h0695: data_out = 8'h8F;
                    16'h0696: data_out = 8'h90;
                    16'h0697: data_out = 8'h91;
                    16'h0698: data_out = 8'h92;
                    16'h0699: data_out = 8'h93;
                    16'h069A: data_out = 8'h94;
                    16'h069B: data_out = 8'h95;
                    16'h069C: data_out = 8'h96;
                    16'h069D: data_out = 8'h97;
                    16'h069E: data_out = 8'h98;
                    16'h069F: data_out = 8'h99;
                    16'h06A0: data_out = 8'h9A;
                    16'h06A1: data_out = 8'h9B;
                    16'h06A2: data_out = 8'h9C;
                    16'h06A3: data_out = 8'h9D;
                    16'h06A4: data_out = 8'h9E;
                    16'h06A5: data_out = 8'h9F;
                    16'h06A6: data_out = 8'hA0;
                    16'h06A7: data_out = 8'hA1;
                    16'h06A8: data_out = 8'hA2;
                    16'h06A9: data_out = 8'hA3;
                    16'h06AA: data_out = 8'hA4;
                    16'h06AB: data_out = 8'hA5;
                    16'h06AC: data_out = 8'hA6;
                    16'h06AD: data_out = 8'hA7;
                    16'h06AE: data_out = 8'hA8;
                    16'h06AF: data_out = 8'hA9;
                    16'h06B0: data_out = 8'hAA;
                    16'h06B1: data_out = 8'hAB;
                    16'h06B2: data_out = 8'hAC;
                    16'h06B3: data_out = 8'hAD;
                    16'h06B4: data_out = 8'hAE;
                    16'h06B5: data_out = 8'hAF;
                    16'h06B6: data_out = 8'hB0;
                    16'h06B7: data_out = 8'hB1;
                    16'h06B8: data_out = 8'hB2;
                    16'h06B9: data_out = 8'hB3;
                    16'h06BA: data_out = 8'hB4;
                    16'h06BB: data_out = 8'hB5;
                    16'h06BC: data_out = 8'hB6;
                    16'h06BD: data_out = 8'hB7;
                    16'h06BE: data_out = 8'hB8;
                    16'h06BF: data_out = 8'hB9;
                    16'h06C0: data_out = 8'hBA;
                    16'h06C1: data_out = 8'hBB;
                    16'h06C2: data_out = 8'hBC;
                    16'h06C3: data_out = 8'hBD;
                    16'h06C4: data_out = 8'hBE;
                    16'h06C5: data_out = 8'hBF;
                    16'h06C6: data_out = 8'hC0;
                    16'h06C7: data_out = 8'hC1;
                    16'h06C8: data_out = 8'hC2;
                    16'h06C9: data_out = 8'hC3;
                    16'h06CA: data_out = 8'hC4;
                    16'h06CB: data_out = 8'hC5;
                    16'h06CC: data_out = 8'hC6;
                    16'h06CD: data_out = 8'hC7;
                    16'h06CE: data_out = 8'hC8;
                    16'h06CF: data_out = 8'hC9;
                    16'h06D0: data_out = 8'hCA;
                    16'h06D1: data_out = 8'hCB;
                    16'h06D2: data_out = 8'hCC;
                    16'h06D3: data_out = 8'hCD;
                    16'h06D4: data_out = 8'hCE;
                    16'h06D5: data_out = 8'hCF;
                    16'h06D6: data_out = 8'hD0;
                    16'h06D7: data_out = 8'hD1;
                    16'h06D8: data_out = 8'hD2;
                    16'h06D9: data_out = 8'hD3;
                    16'h06DA: data_out = 8'hD4;
                    16'h06DB: data_out = 8'hD5;
                    16'h06DC: data_out = 8'hD6;
                    16'h06DD: data_out = 8'hD7;
                    16'h06DE: data_out = 8'hD8;
                    16'h06DF: data_out = 8'hD9;
                    16'h06E0: data_out = 8'hDA;
                    16'h06E1: data_out = 8'hDB;
                    16'h06E2: data_out = 8'hDC;
                    16'h06E3: data_out = 8'hDD;
                    16'h06E4: data_out = 8'hDE;
                    16'h06E5: data_out = 8'hDF;
                    16'h06E6: data_out = 8'hE0;
                    16'h06E7: data_out = 8'hE1;
                    16'h06E8: data_out = 8'hE2;
                    16'h06E9: data_out = 8'hE3;
                    16'h06EA: data_out = 8'hE4;
                    16'h06EB: data_out = 8'hE5;
                    16'h06EC: data_out = 8'hE6;
                    16'h06ED: data_out = 8'hE7;
                    16'h06EE: data_out = 8'hE8;
                    16'h06EF: data_out = 8'hE9;
                    16'h06F0: data_out = 8'hEA;
                    16'h06F1: data_out = 8'hEB;
                    16'h06F2: data_out = 8'hEC;
                    16'h06F3: data_out = 8'hED;
                    16'h06F4: data_out = 8'hEE;
                    16'h06F5: data_out = 8'hEF;
                    16'h06F6: data_out = 8'hF0;
                    16'h06F7: data_out = 8'hF1;
                    16'h06F8: data_out = 8'hF2;
                    16'h06F9: data_out = 8'hF3;
                    16'h06FA: data_out = 8'hF4;
                    16'h06FB: data_out = 8'hF5;
                    16'h06FC: data_out = 8'hF6;
                    16'h06FD: data_out = 8'hF7;
                    16'h06FE: data_out = 8'hF8;
                    16'h06FF: data_out = 8'hF9;
                    16'h0700: data_out = 8'h7;
                    16'h0701: data_out = 8'h8;
                    16'h0702: data_out = 8'h9;
                    16'h0703: data_out = 8'hA;
                    16'h0704: data_out = 8'hB;
                    16'h0705: data_out = 8'hC;
                    16'h0706: data_out = 8'hD;
                    16'h0707: data_out = 8'hE;
                    16'h0708: data_out = 8'hF;
                    16'h0709: data_out = 8'h10;
                    16'h070A: data_out = 8'h11;
                    16'h070B: data_out = 8'h12;
                    16'h070C: data_out = 8'h13;
                    16'h070D: data_out = 8'h14;
                    16'h070E: data_out = 8'h15;
                    16'h070F: data_out = 8'h16;
                    16'h0710: data_out = 8'h17;
                    16'h0711: data_out = 8'h18;
                    16'h0712: data_out = 8'h19;
                    16'h0713: data_out = 8'h1A;
                    16'h0714: data_out = 8'h1B;
                    16'h0715: data_out = 8'h1C;
                    16'h0716: data_out = 8'h1D;
                    16'h0717: data_out = 8'h1E;
                    16'h0718: data_out = 8'h1F;
                    16'h0719: data_out = 8'h20;
                    16'h071A: data_out = 8'h21;
                    16'h071B: data_out = 8'h22;
                    16'h071C: data_out = 8'h23;
                    16'h071D: data_out = 8'h24;
                    16'h071E: data_out = 8'h25;
                    16'h071F: data_out = 8'h26;
                    16'h0720: data_out = 8'h27;
                    16'h0721: data_out = 8'h28;
                    16'h0722: data_out = 8'h29;
                    16'h0723: data_out = 8'h2A;
                    16'h0724: data_out = 8'h2B;
                    16'h0725: data_out = 8'h2C;
                    16'h0726: data_out = 8'h2D;
                    16'h0727: data_out = 8'h2E;
                    16'h0728: data_out = 8'h2F;
                    16'h0729: data_out = 8'h30;
                    16'h072A: data_out = 8'h31;
                    16'h072B: data_out = 8'h32;
                    16'h072C: data_out = 8'h33;
                    16'h072D: data_out = 8'h34;
                    16'h072E: data_out = 8'h35;
                    16'h072F: data_out = 8'h36;
                    16'h0730: data_out = 8'h37;
                    16'h0731: data_out = 8'h38;
                    16'h0732: data_out = 8'h39;
                    16'h0733: data_out = 8'h3A;
                    16'h0734: data_out = 8'h3B;
                    16'h0735: data_out = 8'h3C;
                    16'h0736: data_out = 8'h3D;
                    16'h0737: data_out = 8'h3E;
                    16'h0738: data_out = 8'h3F;
                    16'h0739: data_out = 8'h40;
                    16'h073A: data_out = 8'h41;
                    16'h073B: data_out = 8'h42;
                    16'h073C: data_out = 8'h43;
                    16'h073D: data_out = 8'h44;
                    16'h073E: data_out = 8'h45;
                    16'h073F: data_out = 8'h46;
                    16'h0740: data_out = 8'h47;
                    16'h0741: data_out = 8'h48;
                    16'h0742: data_out = 8'h49;
                    16'h0743: data_out = 8'h4A;
                    16'h0744: data_out = 8'h4B;
                    16'h0745: data_out = 8'h4C;
                    16'h0746: data_out = 8'h4D;
                    16'h0747: data_out = 8'h4E;
                    16'h0748: data_out = 8'h4F;
                    16'h0749: data_out = 8'h50;
                    16'h074A: data_out = 8'h51;
                    16'h074B: data_out = 8'h52;
                    16'h074C: data_out = 8'h53;
                    16'h074D: data_out = 8'h54;
                    16'h074E: data_out = 8'h55;
                    16'h074F: data_out = 8'h56;
                    16'h0750: data_out = 8'h57;
                    16'h0751: data_out = 8'h58;
                    16'h0752: data_out = 8'h59;
                    16'h0753: data_out = 8'h5A;
                    16'h0754: data_out = 8'h5B;
                    16'h0755: data_out = 8'h5C;
                    16'h0756: data_out = 8'h5D;
                    16'h0757: data_out = 8'h5E;
                    16'h0758: data_out = 8'h5F;
                    16'h0759: data_out = 8'h60;
                    16'h075A: data_out = 8'h61;
                    16'h075B: data_out = 8'h62;
                    16'h075C: data_out = 8'h63;
                    16'h075D: data_out = 8'h64;
                    16'h075E: data_out = 8'h65;
                    16'h075F: data_out = 8'h66;
                    16'h0760: data_out = 8'h67;
                    16'h0761: data_out = 8'h68;
                    16'h0762: data_out = 8'h69;
                    16'h0763: data_out = 8'h6A;
                    16'h0764: data_out = 8'h6B;
                    16'h0765: data_out = 8'h6C;
                    16'h0766: data_out = 8'h6D;
                    16'h0767: data_out = 8'h6E;
                    16'h0768: data_out = 8'h6F;
                    16'h0769: data_out = 8'h70;
                    16'h076A: data_out = 8'h71;
                    16'h076B: data_out = 8'h72;
                    16'h076C: data_out = 8'h73;
                    16'h076D: data_out = 8'h74;
                    16'h076E: data_out = 8'h75;
                    16'h076F: data_out = 8'h76;
                    16'h0770: data_out = 8'h77;
                    16'h0771: data_out = 8'h78;
                    16'h0772: data_out = 8'h79;
                    16'h0773: data_out = 8'h7A;
                    16'h0774: data_out = 8'h7B;
                    16'h0775: data_out = 8'h7C;
                    16'h0776: data_out = 8'h7D;
                    16'h0777: data_out = 8'h7E;
                    16'h0778: data_out = 8'h7F;
                    16'h0779: data_out = 8'h80;
                    16'h077A: data_out = 8'h81;
                    16'h077B: data_out = 8'h82;
                    16'h077C: data_out = 8'h83;
                    16'h077D: data_out = 8'h84;
                    16'h077E: data_out = 8'h85;
                    16'h077F: data_out = 8'h86;
                    16'h0780: data_out = 8'h7;
                    16'h0781: data_out = 8'h6;
                    16'h0782: data_out = 8'h5;
                    16'h0783: data_out = 8'h4;
                    16'h0784: data_out = 8'h3;
                    16'h0785: data_out = 8'h2;
                    16'h0786: data_out = 8'h1;
                    16'h0787: data_out = 8'h0;
                    16'h0788: data_out = 8'h81;
                    16'h0789: data_out = 8'h82;
                    16'h078A: data_out = 8'h83;
                    16'h078B: data_out = 8'h84;
                    16'h078C: data_out = 8'h85;
                    16'h078D: data_out = 8'h86;
                    16'h078E: data_out = 8'h87;
                    16'h078F: data_out = 8'h88;
                    16'h0790: data_out = 8'h89;
                    16'h0791: data_out = 8'h8A;
                    16'h0792: data_out = 8'h8B;
                    16'h0793: data_out = 8'h8C;
                    16'h0794: data_out = 8'h8D;
                    16'h0795: data_out = 8'h8E;
                    16'h0796: data_out = 8'h8F;
                    16'h0797: data_out = 8'h90;
                    16'h0798: data_out = 8'h91;
                    16'h0799: data_out = 8'h92;
                    16'h079A: data_out = 8'h93;
                    16'h079B: data_out = 8'h94;
                    16'h079C: data_out = 8'h95;
                    16'h079D: data_out = 8'h96;
                    16'h079E: data_out = 8'h97;
                    16'h079F: data_out = 8'h98;
                    16'h07A0: data_out = 8'h99;
                    16'h07A1: data_out = 8'h9A;
                    16'h07A2: data_out = 8'h9B;
                    16'h07A3: data_out = 8'h9C;
                    16'h07A4: data_out = 8'h9D;
                    16'h07A5: data_out = 8'h9E;
                    16'h07A6: data_out = 8'h9F;
                    16'h07A7: data_out = 8'hA0;
                    16'h07A8: data_out = 8'hA1;
                    16'h07A9: data_out = 8'hA2;
                    16'h07AA: data_out = 8'hA3;
                    16'h07AB: data_out = 8'hA4;
                    16'h07AC: data_out = 8'hA5;
                    16'h07AD: data_out = 8'hA6;
                    16'h07AE: data_out = 8'hA7;
                    16'h07AF: data_out = 8'hA8;
                    16'h07B0: data_out = 8'hA9;
                    16'h07B1: data_out = 8'hAA;
                    16'h07B2: data_out = 8'hAB;
                    16'h07B3: data_out = 8'hAC;
                    16'h07B4: data_out = 8'hAD;
                    16'h07B5: data_out = 8'hAE;
                    16'h07B6: data_out = 8'hAF;
                    16'h07B7: data_out = 8'hB0;
                    16'h07B8: data_out = 8'hB1;
                    16'h07B9: data_out = 8'hB2;
                    16'h07BA: data_out = 8'hB3;
                    16'h07BB: data_out = 8'hB4;
                    16'h07BC: data_out = 8'hB5;
                    16'h07BD: data_out = 8'hB6;
                    16'h07BE: data_out = 8'hB7;
                    16'h07BF: data_out = 8'hB8;
                    16'h07C0: data_out = 8'hB9;
                    16'h07C1: data_out = 8'hBA;
                    16'h07C2: data_out = 8'hBB;
                    16'h07C3: data_out = 8'hBC;
                    16'h07C4: data_out = 8'hBD;
                    16'h07C5: data_out = 8'hBE;
                    16'h07C6: data_out = 8'hBF;
                    16'h07C7: data_out = 8'hC0;
                    16'h07C8: data_out = 8'hC1;
                    16'h07C9: data_out = 8'hC2;
                    16'h07CA: data_out = 8'hC3;
                    16'h07CB: data_out = 8'hC4;
                    16'h07CC: data_out = 8'hC5;
                    16'h07CD: data_out = 8'hC6;
                    16'h07CE: data_out = 8'hC7;
                    16'h07CF: data_out = 8'hC8;
                    16'h07D0: data_out = 8'hC9;
                    16'h07D1: data_out = 8'hCA;
                    16'h07D2: data_out = 8'hCB;
                    16'h07D3: data_out = 8'hCC;
                    16'h07D4: data_out = 8'hCD;
                    16'h07D5: data_out = 8'hCE;
                    16'h07D6: data_out = 8'hCF;
                    16'h07D7: data_out = 8'hD0;
                    16'h07D8: data_out = 8'hD1;
                    16'h07D9: data_out = 8'hD2;
                    16'h07DA: data_out = 8'hD3;
                    16'h07DB: data_out = 8'hD4;
                    16'h07DC: data_out = 8'hD5;
                    16'h07DD: data_out = 8'hD6;
                    16'h07DE: data_out = 8'hD7;
                    16'h07DF: data_out = 8'hD8;
                    16'h07E0: data_out = 8'hD9;
                    16'h07E1: data_out = 8'hDA;
                    16'h07E2: data_out = 8'hDB;
                    16'h07E3: data_out = 8'hDC;
                    16'h07E4: data_out = 8'hDD;
                    16'h07E5: data_out = 8'hDE;
                    16'h07E6: data_out = 8'hDF;
                    16'h07E7: data_out = 8'hE0;
                    16'h07E8: data_out = 8'hE1;
                    16'h07E9: data_out = 8'hE2;
                    16'h07EA: data_out = 8'hE3;
                    16'h07EB: data_out = 8'hE4;
                    16'h07EC: data_out = 8'hE5;
                    16'h07ED: data_out = 8'hE6;
                    16'h07EE: data_out = 8'hE7;
                    16'h07EF: data_out = 8'hE8;
                    16'h07F0: data_out = 8'hE9;
                    16'h07F1: data_out = 8'hEA;
                    16'h07F2: data_out = 8'hEB;
                    16'h07F3: data_out = 8'hEC;
                    16'h07F4: data_out = 8'hED;
                    16'h07F5: data_out = 8'hEE;
                    16'h07F6: data_out = 8'hEF;
                    16'h07F7: data_out = 8'hF0;
                    16'h07F8: data_out = 8'hF1;
                    16'h07F9: data_out = 8'hF2;
                    16'h07FA: data_out = 8'hF3;
                    16'h07FB: data_out = 8'hF4;
                    16'h07FC: data_out = 8'hF5;
                    16'h07FD: data_out = 8'hF6;
                    16'h07FE: data_out = 8'hF7;
                    16'h07FF: data_out = 8'hF8;
                    16'h0800: data_out = 8'h8;
                    16'h0801: data_out = 8'h9;
                    16'h0802: data_out = 8'hA;
                    16'h0803: data_out = 8'hB;
                    16'h0804: data_out = 8'hC;
                    16'h0805: data_out = 8'hD;
                    16'h0806: data_out = 8'hE;
                    16'h0807: data_out = 8'hF;
                    16'h0808: data_out = 8'h10;
                    16'h0809: data_out = 8'h11;
                    16'h080A: data_out = 8'h12;
                    16'h080B: data_out = 8'h13;
                    16'h080C: data_out = 8'h14;
                    16'h080D: data_out = 8'h15;
                    16'h080E: data_out = 8'h16;
                    16'h080F: data_out = 8'h17;
                    16'h0810: data_out = 8'h18;
                    16'h0811: data_out = 8'h19;
                    16'h0812: data_out = 8'h1A;
                    16'h0813: data_out = 8'h1B;
                    16'h0814: data_out = 8'h1C;
                    16'h0815: data_out = 8'h1D;
                    16'h0816: data_out = 8'h1E;
                    16'h0817: data_out = 8'h1F;
                    16'h0818: data_out = 8'h20;
                    16'h0819: data_out = 8'h21;
                    16'h081A: data_out = 8'h22;
                    16'h081B: data_out = 8'h23;
                    16'h081C: data_out = 8'h24;
                    16'h081D: data_out = 8'h25;
                    16'h081E: data_out = 8'h26;
                    16'h081F: data_out = 8'h27;
                    16'h0820: data_out = 8'h28;
                    16'h0821: data_out = 8'h29;
                    16'h0822: data_out = 8'h2A;
                    16'h0823: data_out = 8'h2B;
                    16'h0824: data_out = 8'h2C;
                    16'h0825: data_out = 8'h2D;
                    16'h0826: data_out = 8'h2E;
                    16'h0827: data_out = 8'h2F;
                    16'h0828: data_out = 8'h30;
                    16'h0829: data_out = 8'h31;
                    16'h082A: data_out = 8'h32;
                    16'h082B: data_out = 8'h33;
                    16'h082C: data_out = 8'h34;
                    16'h082D: data_out = 8'h35;
                    16'h082E: data_out = 8'h36;
                    16'h082F: data_out = 8'h37;
                    16'h0830: data_out = 8'h38;
                    16'h0831: data_out = 8'h39;
                    16'h0832: data_out = 8'h3A;
                    16'h0833: data_out = 8'h3B;
                    16'h0834: data_out = 8'h3C;
                    16'h0835: data_out = 8'h3D;
                    16'h0836: data_out = 8'h3E;
                    16'h0837: data_out = 8'h3F;
                    16'h0838: data_out = 8'h40;
                    16'h0839: data_out = 8'h41;
                    16'h083A: data_out = 8'h42;
                    16'h083B: data_out = 8'h43;
                    16'h083C: data_out = 8'h44;
                    16'h083D: data_out = 8'h45;
                    16'h083E: data_out = 8'h46;
                    16'h083F: data_out = 8'h47;
                    16'h0840: data_out = 8'h48;
                    16'h0841: data_out = 8'h49;
                    16'h0842: data_out = 8'h4A;
                    16'h0843: data_out = 8'h4B;
                    16'h0844: data_out = 8'h4C;
                    16'h0845: data_out = 8'h4D;
                    16'h0846: data_out = 8'h4E;
                    16'h0847: data_out = 8'h4F;
                    16'h0848: data_out = 8'h50;
                    16'h0849: data_out = 8'h51;
                    16'h084A: data_out = 8'h52;
                    16'h084B: data_out = 8'h53;
                    16'h084C: data_out = 8'h54;
                    16'h084D: data_out = 8'h55;
                    16'h084E: data_out = 8'h56;
                    16'h084F: data_out = 8'h57;
                    16'h0850: data_out = 8'h58;
                    16'h0851: data_out = 8'h59;
                    16'h0852: data_out = 8'h5A;
                    16'h0853: data_out = 8'h5B;
                    16'h0854: data_out = 8'h5C;
                    16'h0855: data_out = 8'h5D;
                    16'h0856: data_out = 8'h5E;
                    16'h0857: data_out = 8'h5F;
                    16'h0858: data_out = 8'h60;
                    16'h0859: data_out = 8'h61;
                    16'h085A: data_out = 8'h62;
                    16'h085B: data_out = 8'h63;
                    16'h085C: data_out = 8'h64;
                    16'h085D: data_out = 8'h65;
                    16'h085E: data_out = 8'h66;
                    16'h085F: data_out = 8'h67;
                    16'h0860: data_out = 8'h68;
                    16'h0861: data_out = 8'h69;
                    16'h0862: data_out = 8'h6A;
                    16'h0863: data_out = 8'h6B;
                    16'h0864: data_out = 8'h6C;
                    16'h0865: data_out = 8'h6D;
                    16'h0866: data_out = 8'h6E;
                    16'h0867: data_out = 8'h6F;
                    16'h0868: data_out = 8'h70;
                    16'h0869: data_out = 8'h71;
                    16'h086A: data_out = 8'h72;
                    16'h086B: data_out = 8'h73;
                    16'h086C: data_out = 8'h74;
                    16'h086D: data_out = 8'h75;
                    16'h086E: data_out = 8'h76;
                    16'h086F: data_out = 8'h77;
                    16'h0870: data_out = 8'h78;
                    16'h0871: data_out = 8'h79;
                    16'h0872: data_out = 8'h7A;
                    16'h0873: data_out = 8'h7B;
                    16'h0874: data_out = 8'h7C;
                    16'h0875: data_out = 8'h7D;
                    16'h0876: data_out = 8'h7E;
                    16'h0877: data_out = 8'h7F;
                    16'h0878: data_out = 8'h80;
                    16'h0879: data_out = 8'h81;
                    16'h087A: data_out = 8'h82;
                    16'h087B: data_out = 8'h83;
                    16'h087C: data_out = 8'h84;
                    16'h087D: data_out = 8'h85;
                    16'h087E: data_out = 8'h86;
                    16'h087F: data_out = 8'h87;
                    16'h0880: data_out = 8'h8;
                    16'h0881: data_out = 8'h7;
                    16'h0882: data_out = 8'h6;
                    16'h0883: data_out = 8'h5;
                    16'h0884: data_out = 8'h4;
                    16'h0885: data_out = 8'h3;
                    16'h0886: data_out = 8'h2;
                    16'h0887: data_out = 8'h1;
                    16'h0888: data_out = 8'h0;
                    16'h0889: data_out = 8'h81;
                    16'h088A: data_out = 8'h82;
                    16'h088B: data_out = 8'h83;
                    16'h088C: data_out = 8'h84;
                    16'h088D: data_out = 8'h85;
                    16'h088E: data_out = 8'h86;
                    16'h088F: data_out = 8'h87;
                    16'h0890: data_out = 8'h88;
                    16'h0891: data_out = 8'h89;
                    16'h0892: data_out = 8'h8A;
                    16'h0893: data_out = 8'h8B;
                    16'h0894: data_out = 8'h8C;
                    16'h0895: data_out = 8'h8D;
                    16'h0896: data_out = 8'h8E;
                    16'h0897: data_out = 8'h8F;
                    16'h0898: data_out = 8'h90;
                    16'h0899: data_out = 8'h91;
                    16'h089A: data_out = 8'h92;
                    16'h089B: data_out = 8'h93;
                    16'h089C: data_out = 8'h94;
                    16'h089D: data_out = 8'h95;
                    16'h089E: data_out = 8'h96;
                    16'h089F: data_out = 8'h97;
                    16'h08A0: data_out = 8'h98;
                    16'h08A1: data_out = 8'h99;
                    16'h08A2: data_out = 8'h9A;
                    16'h08A3: data_out = 8'h9B;
                    16'h08A4: data_out = 8'h9C;
                    16'h08A5: data_out = 8'h9D;
                    16'h08A6: data_out = 8'h9E;
                    16'h08A7: data_out = 8'h9F;
                    16'h08A8: data_out = 8'hA0;
                    16'h08A9: data_out = 8'hA1;
                    16'h08AA: data_out = 8'hA2;
                    16'h08AB: data_out = 8'hA3;
                    16'h08AC: data_out = 8'hA4;
                    16'h08AD: data_out = 8'hA5;
                    16'h08AE: data_out = 8'hA6;
                    16'h08AF: data_out = 8'hA7;
                    16'h08B0: data_out = 8'hA8;
                    16'h08B1: data_out = 8'hA9;
                    16'h08B2: data_out = 8'hAA;
                    16'h08B3: data_out = 8'hAB;
                    16'h08B4: data_out = 8'hAC;
                    16'h08B5: data_out = 8'hAD;
                    16'h08B6: data_out = 8'hAE;
                    16'h08B7: data_out = 8'hAF;
                    16'h08B8: data_out = 8'hB0;
                    16'h08B9: data_out = 8'hB1;
                    16'h08BA: data_out = 8'hB2;
                    16'h08BB: data_out = 8'hB3;
                    16'h08BC: data_out = 8'hB4;
                    16'h08BD: data_out = 8'hB5;
                    16'h08BE: data_out = 8'hB6;
                    16'h08BF: data_out = 8'hB7;
                    16'h08C0: data_out = 8'hB8;
                    16'h08C1: data_out = 8'hB9;
                    16'h08C2: data_out = 8'hBA;
                    16'h08C3: data_out = 8'hBB;
                    16'h08C4: data_out = 8'hBC;
                    16'h08C5: data_out = 8'hBD;
                    16'h08C6: data_out = 8'hBE;
                    16'h08C7: data_out = 8'hBF;
                    16'h08C8: data_out = 8'hC0;
                    16'h08C9: data_out = 8'hC1;
                    16'h08CA: data_out = 8'hC2;
                    16'h08CB: data_out = 8'hC3;
                    16'h08CC: data_out = 8'hC4;
                    16'h08CD: data_out = 8'hC5;
                    16'h08CE: data_out = 8'hC6;
                    16'h08CF: data_out = 8'hC7;
                    16'h08D0: data_out = 8'hC8;
                    16'h08D1: data_out = 8'hC9;
                    16'h08D2: data_out = 8'hCA;
                    16'h08D3: data_out = 8'hCB;
                    16'h08D4: data_out = 8'hCC;
                    16'h08D5: data_out = 8'hCD;
                    16'h08D6: data_out = 8'hCE;
                    16'h08D7: data_out = 8'hCF;
                    16'h08D8: data_out = 8'hD0;
                    16'h08D9: data_out = 8'hD1;
                    16'h08DA: data_out = 8'hD2;
                    16'h08DB: data_out = 8'hD3;
                    16'h08DC: data_out = 8'hD4;
                    16'h08DD: data_out = 8'hD5;
                    16'h08DE: data_out = 8'hD6;
                    16'h08DF: data_out = 8'hD7;
                    16'h08E0: data_out = 8'hD8;
                    16'h08E1: data_out = 8'hD9;
                    16'h08E2: data_out = 8'hDA;
                    16'h08E3: data_out = 8'hDB;
                    16'h08E4: data_out = 8'hDC;
                    16'h08E5: data_out = 8'hDD;
                    16'h08E6: data_out = 8'hDE;
                    16'h08E7: data_out = 8'hDF;
                    16'h08E8: data_out = 8'hE0;
                    16'h08E9: data_out = 8'hE1;
                    16'h08EA: data_out = 8'hE2;
                    16'h08EB: data_out = 8'hE3;
                    16'h08EC: data_out = 8'hE4;
                    16'h08ED: data_out = 8'hE5;
                    16'h08EE: data_out = 8'hE6;
                    16'h08EF: data_out = 8'hE7;
                    16'h08F0: data_out = 8'hE8;
                    16'h08F1: data_out = 8'hE9;
                    16'h08F2: data_out = 8'hEA;
                    16'h08F3: data_out = 8'hEB;
                    16'h08F4: data_out = 8'hEC;
                    16'h08F5: data_out = 8'hED;
                    16'h08F6: data_out = 8'hEE;
                    16'h08F7: data_out = 8'hEF;
                    16'h08F8: data_out = 8'hF0;
                    16'h08F9: data_out = 8'hF1;
                    16'h08FA: data_out = 8'hF2;
                    16'h08FB: data_out = 8'hF3;
                    16'h08FC: data_out = 8'hF4;
                    16'h08FD: data_out = 8'hF5;
                    16'h08FE: data_out = 8'hF6;
                    16'h08FF: data_out = 8'hF7;
                    16'h0900: data_out = 8'h9;
                    16'h0901: data_out = 8'hA;
                    16'h0902: data_out = 8'hB;
                    16'h0903: data_out = 8'hC;
                    16'h0904: data_out = 8'hD;
                    16'h0905: data_out = 8'hE;
                    16'h0906: data_out = 8'hF;
                    16'h0907: data_out = 8'h10;
                    16'h0908: data_out = 8'h11;
                    16'h0909: data_out = 8'h12;
                    16'h090A: data_out = 8'h13;
                    16'h090B: data_out = 8'h14;
                    16'h090C: data_out = 8'h15;
                    16'h090D: data_out = 8'h16;
                    16'h090E: data_out = 8'h17;
                    16'h090F: data_out = 8'h18;
                    16'h0910: data_out = 8'h19;
                    16'h0911: data_out = 8'h1A;
                    16'h0912: data_out = 8'h1B;
                    16'h0913: data_out = 8'h1C;
                    16'h0914: data_out = 8'h1D;
                    16'h0915: data_out = 8'h1E;
                    16'h0916: data_out = 8'h1F;
                    16'h0917: data_out = 8'h20;
                    16'h0918: data_out = 8'h21;
                    16'h0919: data_out = 8'h22;
                    16'h091A: data_out = 8'h23;
                    16'h091B: data_out = 8'h24;
                    16'h091C: data_out = 8'h25;
                    16'h091D: data_out = 8'h26;
                    16'h091E: data_out = 8'h27;
                    16'h091F: data_out = 8'h28;
                    16'h0920: data_out = 8'h29;
                    16'h0921: data_out = 8'h2A;
                    16'h0922: data_out = 8'h2B;
                    16'h0923: data_out = 8'h2C;
                    16'h0924: data_out = 8'h2D;
                    16'h0925: data_out = 8'h2E;
                    16'h0926: data_out = 8'h2F;
                    16'h0927: data_out = 8'h30;
                    16'h0928: data_out = 8'h31;
                    16'h0929: data_out = 8'h32;
                    16'h092A: data_out = 8'h33;
                    16'h092B: data_out = 8'h34;
                    16'h092C: data_out = 8'h35;
                    16'h092D: data_out = 8'h36;
                    16'h092E: data_out = 8'h37;
                    16'h092F: data_out = 8'h38;
                    16'h0930: data_out = 8'h39;
                    16'h0931: data_out = 8'h3A;
                    16'h0932: data_out = 8'h3B;
                    16'h0933: data_out = 8'h3C;
                    16'h0934: data_out = 8'h3D;
                    16'h0935: data_out = 8'h3E;
                    16'h0936: data_out = 8'h3F;
                    16'h0937: data_out = 8'h40;
                    16'h0938: data_out = 8'h41;
                    16'h0939: data_out = 8'h42;
                    16'h093A: data_out = 8'h43;
                    16'h093B: data_out = 8'h44;
                    16'h093C: data_out = 8'h45;
                    16'h093D: data_out = 8'h46;
                    16'h093E: data_out = 8'h47;
                    16'h093F: data_out = 8'h48;
                    16'h0940: data_out = 8'h49;
                    16'h0941: data_out = 8'h4A;
                    16'h0942: data_out = 8'h4B;
                    16'h0943: data_out = 8'h4C;
                    16'h0944: data_out = 8'h4D;
                    16'h0945: data_out = 8'h4E;
                    16'h0946: data_out = 8'h4F;
                    16'h0947: data_out = 8'h50;
                    16'h0948: data_out = 8'h51;
                    16'h0949: data_out = 8'h52;
                    16'h094A: data_out = 8'h53;
                    16'h094B: data_out = 8'h54;
                    16'h094C: data_out = 8'h55;
                    16'h094D: data_out = 8'h56;
                    16'h094E: data_out = 8'h57;
                    16'h094F: data_out = 8'h58;
                    16'h0950: data_out = 8'h59;
                    16'h0951: data_out = 8'h5A;
                    16'h0952: data_out = 8'h5B;
                    16'h0953: data_out = 8'h5C;
                    16'h0954: data_out = 8'h5D;
                    16'h0955: data_out = 8'h5E;
                    16'h0956: data_out = 8'h5F;
                    16'h0957: data_out = 8'h60;
                    16'h0958: data_out = 8'h61;
                    16'h0959: data_out = 8'h62;
                    16'h095A: data_out = 8'h63;
                    16'h095B: data_out = 8'h64;
                    16'h095C: data_out = 8'h65;
                    16'h095D: data_out = 8'h66;
                    16'h095E: data_out = 8'h67;
                    16'h095F: data_out = 8'h68;
                    16'h0960: data_out = 8'h69;
                    16'h0961: data_out = 8'h6A;
                    16'h0962: data_out = 8'h6B;
                    16'h0963: data_out = 8'h6C;
                    16'h0964: data_out = 8'h6D;
                    16'h0965: data_out = 8'h6E;
                    16'h0966: data_out = 8'h6F;
                    16'h0967: data_out = 8'h70;
                    16'h0968: data_out = 8'h71;
                    16'h0969: data_out = 8'h72;
                    16'h096A: data_out = 8'h73;
                    16'h096B: data_out = 8'h74;
                    16'h096C: data_out = 8'h75;
                    16'h096D: data_out = 8'h76;
                    16'h096E: data_out = 8'h77;
                    16'h096F: data_out = 8'h78;
                    16'h0970: data_out = 8'h79;
                    16'h0971: data_out = 8'h7A;
                    16'h0972: data_out = 8'h7B;
                    16'h0973: data_out = 8'h7C;
                    16'h0974: data_out = 8'h7D;
                    16'h0975: data_out = 8'h7E;
                    16'h0976: data_out = 8'h7F;
                    16'h0977: data_out = 8'h80;
                    16'h0978: data_out = 8'h81;
                    16'h0979: data_out = 8'h82;
                    16'h097A: data_out = 8'h83;
                    16'h097B: data_out = 8'h84;
                    16'h097C: data_out = 8'h85;
                    16'h097D: data_out = 8'h86;
                    16'h097E: data_out = 8'h87;
                    16'h097F: data_out = 8'h88;
                    16'h0980: data_out = 8'h9;
                    16'h0981: data_out = 8'h8;
                    16'h0982: data_out = 8'h7;
                    16'h0983: data_out = 8'h6;
                    16'h0984: data_out = 8'h5;
                    16'h0985: data_out = 8'h4;
                    16'h0986: data_out = 8'h3;
                    16'h0987: data_out = 8'h2;
                    16'h0988: data_out = 8'h1;
                    16'h0989: data_out = 8'h0;
                    16'h098A: data_out = 8'h81;
                    16'h098B: data_out = 8'h82;
                    16'h098C: data_out = 8'h83;
                    16'h098D: data_out = 8'h84;
                    16'h098E: data_out = 8'h85;
                    16'h098F: data_out = 8'h86;
                    16'h0990: data_out = 8'h87;
                    16'h0991: data_out = 8'h88;
                    16'h0992: data_out = 8'h89;
                    16'h0993: data_out = 8'h8A;
                    16'h0994: data_out = 8'h8B;
                    16'h0995: data_out = 8'h8C;
                    16'h0996: data_out = 8'h8D;
                    16'h0997: data_out = 8'h8E;
                    16'h0998: data_out = 8'h8F;
                    16'h0999: data_out = 8'h90;
                    16'h099A: data_out = 8'h91;
                    16'h099B: data_out = 8'h92;
                    16'h099C: data_out = 8'h93;
                    16'h099D: data_out = 8'h94;
                    16'h099E: data_out = 8'h95;
                    16'h099F: data_out = 8'h96;
                    16'h09A0: data_out = 8'h97;
                    16'h09A1: data_out = 8'h98;
                    16'h09A2: data_out = 8'h99;
                    16'h09A3: data_out = 8'h9A;
                    16'h09A4: data_out = 8'h9B;
                    16'h09A5: data_out = 8'h9C;
                    16'h09A6: data_out = 8'h9D;
                    16'h09A7: data_out = 8'h9E;
                    16'h09A8: data_out = 8'h9F;
                    16'h09A9: data_out = 8'hA0;
                    16'h09AA: data_out = 8'hA1;
                    16'h09AB: data_out = 8'hA2;
                    16'h09AC: data_out = 8'hA3;
                    16'h09AD: data_out = 8'hA4;
                    16'h09AE: data_out = 8'hA5;
                    16'h09AF: data_out = 8'hA6;
                    16'h09B0: data_out = 8'hA7;
                    16'h09B1: data_out = 8'hA8;
                    16'h09B2: data_out = 8'hA9;
                    16'h09B3: data_out = 8'hAA;
                    16'h09B4: data_out = 8'hAB;
                    16'h09B5: data_out = 8'hAC;
                    16'h09B6: data_out = 8'hAD;
                    16'h09B7: data_out = 8'hAE;
                    16'h09B8: data_out = 8'hAF;
                    16'h09B9: data_out = 8'hB0;
                    16'h09BA: data_out = 8'hB1;
                    16'h09BB: data_out = 8'hB2;
                    16'h09BC: data_out = 8'hB3;
                    16'h09BD: data_out = 8'hB4;
                    16'h09BE: data_out = 8'hB5;
                    16'h09BF: data_out = 8'hB6;
                    16'h09C0: data_out = 8'hB7;
                    16'h09C1: data_out = 8'hB8;
                    16'h09C2: data_out = 8'hB9;
                    16'h09C3: data_out = 8'hBA;
                    16'h09C4: data_out = 8'hBB;
                    16'h09C5: data_out = 8'hBC;
                    16'h09C6: data_out = 8'hBD;
                    16'h09C7: data_out = 8'hBE;
                    16'h09C8: data_out = 8'hBF;
                    16'h09C9: data_out = 8'hC0;
                    16'h09CA: data_out = 8'hC1;
                    16'h09CB: data_out = 8'hC2;
                    16'h09CC: data_out = 8'hC3;
                    16'h09CD: data_out = 8'hC4;
                    16'h09CE: data_out = 8'hC5;
                    16'h09CF: data_out = 8'hC6;
                    16'h09D0: data_out = 8'hC7;
                    16'h09D1: data_out = 8'hC8;
                    16'h09D2: data_out = 8'hC9;
                    16'h09D3: data_out = 8'hCA;
                    16'h09D4: data_out = 8'hCB;
                    16'h09D5: data_out = 8'hCC;
                    16'h09D6: data_out = 8'hCD;
                    16'h09D7: data_out = 8'hCE;
                    16'h09D8: data_out = 8'hCF;
                    16'h09D9: data_out = 8'hD0;
                    16'h09DA: data_out = 8'hD1;
                    16'h09DB: data_out = 8'hD2;
                    16'h09DC: data_out = 8'hD3;
                    16'h09DD: data_out = 8'hD4;
                    16'h09DE: data_out = 8'hD5;
                    16'h09DF: data_out = 8'hD6;
                    16'h09E0: data_out = 8'hD7;
                    16'h09E1: data_out = 8'hD8;
                    16'h09E2: data_out = 8'hD9;
                    16'h09E3: data_out = 8'hDA;
                    16'h09E4: data_out = 8'hDB;
                    16'h09E5: data_out = 8'hDC;
                    16'h09E6: data_out = 8'hDD;
                    16'h09E7: data_out = 8'hDE;
                    16'h09E8: data_out = 8'hDF;
                    16'h09E9: data_out = 8'hE0;
                    16'h09EA: data_out = 8'hE1;
                    16'h09EB: data_out = 8'hE2;
                    16'h09EC: data_out = 8'hE3;
                    16'h09ED: data_out = 8'hE4;
                    16'h09EE: data_out = 8'hE5;
                    16'h09EF: data_out = 8'hE6;
                    16'h09F0: data_out = 8'hE7;
                    16'h09F1: data_out = 8'hE8;
                    16'h09F2: data_out = 8'hE9;
                    16'h09F3: data_out = 8'hEA;
                    16'h09F4: data_out = 8'hEB;
                    16'h09F5: data_out = 8'hEC;
                    16'h09F6: data_out = 8'hED;
                    16'h09F7: data_out = 8'hEE;
                    16'h09F8: data_out = 8'hEF;
                    16'h09F9: data_out = 8'hF0;
                    16'h09FA: data_out = 8'hF1;
                    16'h09FB: data_out = 8'hF2;
                    16'h09FC: data_out = 8'hF3;
                    16'h09FD: data_out = 8'hF4;
                    16'h09FE: data_out = 8'hF5;
                    16'h09FF: data_out = 8'hF6;
                    16'h0A00: data_out = 8'hA;
                    16'h0A01: data_out = 8'hB;
                    16'h0A02: data_out = 8'hC;
                    16'h0A03: data_out = 8'hD;
                    16'h0A04: data_out = 8'hE;
                    16'h0A05: data_out = 8'hF;
                    16'h0A06: data_out = 8'h10;
                    16'h0A07: data_out = 8'h11;
                    16'h0A08: data_out = 8'h12;
                    16'h0A09: data_out = 8'h13;
                    16'h0A0A: data_out = 8'h14;
                    16'h0A0B: data_out = 8'h15;
                    16'h0A0C: data_out = 8'h16;
                    16'h0A0D: data_out = 8'h17;
                    16'h0A0E: data_out = 8'h18;
                    16'h0A0F: data_out = 8'h19;
                    16'h0A10: data_out = 8'h1A;
                    16'h0A11: data_out = 8'h1B;
                    16'h0A12: data_out = 8'h1C;
                    16'h0A13: data_out = 8'h1D;
                    16'h0A14: data_out = 8'h1E;
                    16'h0A15: data_out = 8'h1F;
                    16'h0A16: data_out = 8'h20;
                    16'h0A17: data_out = 8'h21;
                    16'h0A18: data_out = 8'h22;
                    16'h0A19: data_out = 8'h23;
                    16'h0A1A: data_out = 8'h24;
                    16'h0A1B: data_out = 8'h25;
                    16'h0A1C: data_out = 8'h26;
                    16'h0A1D: data_out = 8'h27;
                    16'h0A1E: data_out = 8'h28;
                    16'h0A1F: data_out = 8'h29;
                    16'h0A20: data_out = 8'h2A;
                    16'h0A21: data_out = 8'h2B;
                    16'h0A22: data_out = 8'h2C;
                    16'h0A23: data_out = 8'h2D;
                    16'h0A24: data_out = 8'h2E;
                    16'h0A25: data_out = 8'h2F;
                    16'h0A26: data_out = 8'h30;
                    16'h0A27: data_out = 8'h31;
                    16'h0A28: data_out = 8'h32;
                    16'h0A29: data_out = 8'h33;
                    16'h0A2A: data_out = 8'h34;
                    16'h0A2B: data_out = 8'h35;
                    16'h0A2C: data_out = 8'h36;
                    16'h0A2D: data_out = 8'h37;
                    16'h0A2E: data_out = 8'h38;
                    16'h0A2F: data_out = 8'h39;
                    16'h0A30: data_out = 8'h3A;
                    16'h0A31: data_out = 8'h3B;
                    16'h0A32: data_out = 8'h3C;
                    16'h0A33: data_out = 8'h3D;
                    16'h0A34: data_out = 8'h3E;
                    16'h0A35: data_out = 8'h3F;
                    16'h0A36: data_out = 8'h40;
                    16'h0A37: data_out = 8'h41;
                    16'h0A38: data_out = 8'h42;
                    16'h0A39: data_out = 8'h43;
                    16'h0A3A: data_out = 8'h44;
                    16'h0A3B: data_out = 8'h45;
                    16'h0A3C: data_out = 8'h46;
                    16'h0A3D: data_out = 8'h47;
                    16'h0A3E: data_out = 8'h48;
                    16'h0A3F: data_out = 8'h49;
                    16'h0A40: data_out = 8'h4A;
                    16'h0A41: data_out = 8'h4B;
                    16'h0A42: data_out = 8'h4C;
                    16'h0A43: data_out = 8'h4D;
                    16'h0A44: data_out = 8'h4E;
                    16'h0A45: data_out = 8'h4F;
                    16'h0A46: data_out = 8'h50;
                    16'h0A47: data_out = 8'h51;
                    16'h0A48: data_out = 8'h52;
                    16'h0A49: data_out = 8'h53;
                    16'h0A4A: data_out = 8'h54;
                    16'h0A4B: data_out = 8'h55;
                    16'h0A4C: data_out = 8'h56;
                    16'h0A4D: data_out = 8'h57;
                    16'h0A4E: data_out = 8'h58;
                    16'h0A4F: data_out = 8'h59;
                    16'h0A50: data_out = 8'h5A;
                    16'h0A51: data_out = 8'h5B;
                    16'h0A52: data_out = 8'h5C;
                    16'h0A53: data_out = 8'h5D;
                    16'h0A54: data_out = 8'h5E;
                    16'h0A55: data_out = 8'h5F;
                    16'h0A56: data_out = 8'h60;
                    16'h0A57: data_out = 8'h61;
                    16'h0A58: data_out = 8'h62;
                    16'h0A59: data_out = 8'h63;
                    16'h0A5A: data_out = 8'h64;
                    16'h0A5B: data_out = 8'h65;
                    16'h0A5C: data_out = 8'h66;
                    16'h0A5D: data_out = 8'h67;
                    16'h0A5E: data_out = 8'h68;
                    16'h0A5F: data_out = 8'h69;
                    16'h0A60: data_out = 8'h6A;
                    16'h0A61: data_out = 8'h6B;
                    16'h0A62: data_out = 8'h6C;
                    16'h0A63: data_out = 8'h6D;
                    16'h0A64: data_out = 8'h6E;
                    16'h0A65: data_out = 8'h6F;
                    16'h0A66: data_out = 8'h70;
                    16'h0A67: data_out = 8'h71;
                    16'h0A68: data_out = 8'h72;
                    16'h0A69: data_out = 8'h73;
                    16'h0A6A: data_out = 8'h74;
                    16'h0A6B: data_out = 8'h75;
                    16'h0A6C: data_out = 8'h76;
                    16'h0A6D: data_out = 8'h77;
                    16'h0A6E: data_out = 8'h78;
                    16'h0A6F: data_out = 8'h79;
                    16'h0A70: data_out = 8'h7A;
                    16'h0A71: data_out = 8'h7B;
                    16'h0A72: data_out = 8'h7C;
                    16'h0A73: data_out = 8'h7D;
                    16'h0A74: data_out = 8'h7E;
                    16'h0A75: data_out = 8'h7F;
                    16'h0A76: data_out = 8'h80;
                    16'h0A77: data_out = 8'h81;
                    16'h0A78: data_out = 8'h82;
                    16'h0A79: data_out = 8'h83;
                    16'h0A7A: data_out = 8'h84;
                    16'h0A7B: data_out = 8'h85;
                    16'h0A7C: data_out = 8'h86;
                    16'h0A7D: data_out = 8'h87;
                    16'h0A7E: data_out = 8'h88;
                    16'h0A7F: data_out = 8'h89;
                    16'h0A80: data_out = 8'hA;
                    16'h0A81: data_out = 8'h9;
                    16'h0A82: data_out = 8'h8;
                    16'h0A83: data_out = 8'h7;
                    16'h0A84: data_out = 8'h6;
                    16'h0A85: data_out = 8'h5;
                    16'h0A86: data_out = 8'h4;
                    16'h0A87: data_out = 8'h3;
                    16'h0A88: data_out = 8'h2;
                    16'h0A89: data_out = 8'h1;
                    16'h0A8A: data_out = 8'h0;
                    16'h0A8B: data_out = 8'h81;
                    16'h0A8C: data_out = 8'h82;
                    16'h0A8D: data_out = 8'h83;
                    16'h0A8E: data_out = 8'h84;
                    16'h0A8F: data_out = 8'h85;
                    16'h0A90: data_out = 8'h86;
                    16'h0A91: data_out = 8'h87;
                    16'h0A92: data_out = 8'h88;
                    16'h0A93: data_out = 8'h89;
                    16'h0A94: data_out = 8'h8A;
                    16'h0A95: data_out = 8'h8B;
                    16'h0A96: data_out = 8'h8C;
                    16'h0A97: data_out = 8'h8D;
                    16'h0A98: data_out = 8'h8E;
                    16'h0A99: data_out = 8'h8F;
                    16'h0A9A: data_out = 8'h90;
                    16'h0A9B: data_out = 8'h91;
                    16'h0A9C: data_out = 8'h92;
                    16'h0A9D: data_out = 8'h93;
                    16'h0A9E: data_out = 8'h94;
                    16'h0A9F: data_out = 8'h95;
                    16'h0AA0: data_out = 8'h96;
                    16'h0AA1: data_out = 8'h97;
                    16'h0AA2: data_out = 8'h98;
                    16'h0AA3: data_out = 8'h99;
                    16'h0AA4: data_out = 8'h9A;
                    16'h0AA5: data_out = 8'h9B;
                    16'h0AA6: data_out = 8'h9C;
                    16'h0AA7: data_out = 8'h9D;
                    16'h0AA8: data_out = 8'h9E;
                    16'h0AA9: data_out = 8'h9F;
                    16'h0AAA: data_out = 8'hA0;
                    16'h0AAB: data_out = 8'hA1;
                    16'h0AAC: data_out = 8'hA2;
                    16'h0AAD: data_out = 8'hA3;
                    16'h0AAE: data_out = 8'hA4;
                    16'h0AAF: data_out = 8'hA5;
                    16'h0AB0: data_out = 8'hA6;
                    16'h0AB1: data_out = 8'hA7;
                    16'h0AB2: data_out = 8'hA8;
                    16'h0AB3: data_out = 8'hA9;
                    16'h0AB4: data_out = 8'hAA;
                    16'h0AB5: data_out = 8'hAB;
                    16'h0AB6: data_out = 8'hAC;
                    16'h0AB7: data_out = 8'hAD;
                    16'h0AB8: data_out = 8'hAE;
                    16'h0AB9: data_out = 8'hAF;
                    16'h0ABA: data_out = 8'hB0;
                    16'h0ABB: data_out = 8'hB1;
                    16'h0ABC: data_out = 8'hB2;
                    16'h0ABD: data_out = 8'hB3;
                    16'h0ABE: data_out = 8'hB4;
                    16'h0ABF: data_out = 8'hB5;
                    16'h0AC0: data_out = 8'hB6;
                    16'h0AC1: data_out = 8'hB7;
                    16'h0AC2: data_out = 8'hB8;
                    16'h0AC3: data_out = 8'hB9;
                    16'h0AC4: data_out = 8'hBA;
                    16'h0AC5: data_out = 8'hBB;
                    16'h0AC6: data_out = 8'hBC;
                    16'h0AC7: data_out = 8'hBD;
                    16'h0AC8: data_out = 8'hBE;
                    16'h0AC9: data_out = 8'hBF;
                    16'h0ACA: data_out = 8'hC0;
                    16'h0ACB: data_out = 8'hC1;
                    16'h0ACC: data_out = 8'hC2;
                    16'h0ACD: data_out = 8'hC3;
                    16'h0ACE: data_out = 8'hC4;
                    16'h0ACF: data_out = 8'hC5;
                    16'h0AD0: data_out = 8'hC6;
                    16'h0AD1: data_out = 8'hC7;
                    16'h0AD2: data_out = 8'hC8;
                    16'h0AD3: data_out = 8'hC9;
                    16'h0AD4: data_out = 8'hCA;
                    16'h0AD5: data_out = 8'hCB;
                    16'h0AD6: data_out = 8'hCC;
                    16'h0AD7: data_out = 8'hCD;
                    16'h0AD8: data_out = 8'hCE;
                    16'h0AD9: data_out = 8'hCF;
                    16'h0ADA: data_out = 8'hD0;
                    16'h0ADB: data_out = 8'hD1;
                    16'h0ADC: data_out = 8'hD2;
                    16'h0ADD: data_out = 8'hD3;
                    16'h0ADE: data_out = 8'hD4;
                    16'h0ADF: data_out = 8'hD5;
                    16'h0AE0: data_out = 8'hD6;
                    16'h0AE1: data_out = 8'hD7;
                    16'h0AE2: data_out = 8'hD8;
                    16'h0AE3: data_out = 8'hD9;
                    16'h0AE4: data_out = 8'hDA;
                    16'h0AE5: data_out = 8'hDB;
                    16'h0AE6: data_out = 8'hDC;
                    16'h0AE7: data_out = 8'hDD;
                    16'h0AE8: data_out = 8'hDE;
                    16'h0AE9: data_out = 8'hDF;
                    16'h0AEA: data_out = 8'hE0;
                    16'h0AEB: data_out = 8'hE1;
                    16'h0AEC: data_out = 8'hE2;
                    16'h0AED: data_out = 8'hE3;
                    16'h0AEE: data_out = 8'hE4;
                    16'h0AEF: data_out = 8'hE5;
                    16'h0AF0: data_out = 8'hE6;
                    16'h0AF1: data_out = 8'hE7;
                    16'h0AF2: data_out = 8'hE8;
                    16'h0AF3: data_out = 8'hE9;
                    16'h0AF4: data_out = 8'hEA;
                    16'h0AF5: data_out = 8'hEB;
                    16'h0AF6: data_out = 8'hEC;
                    16'h0AF7: data_out = 8'hED;
                    16'h0AF8: data_out = 8'hEE;
                    16'h0AF9: data_out = 8'hEF;
                    16'h0AFA: data_out = 8'hF0;
                    16'h0AFB: data_out = 8'hF1;
                    16'h0AFC: data_out = 8'hF2;
                    16'h0AFD: data_out = 8'hF3;
                    16'h0AFE: data_out = 8'hF4;
                    16'h0AFF: data_out = 8'hF5;
                    16'h0B00: data_out = 8'hB;
                    16'h0B01: data_out = 8'hC;
                    16'h0B02: data_out = 8'hD;
                    16'h0B03: data_out = 8'hE;
                    16'h0B04: data_out = 8'hF;
                    16'h0B05: data_out = 8'h10;
                    16'h0B06: data_out = 8'h11;
                    16'h0B07: data_out = 8'h12;
                    16'h0B08: data_out = 8'h13;
                    16'h0B09: data_out = 8'h14;
                    16'h0B0A: data_out = 8'h15;
                    16'h0B0B: data_out = 8'h16;
                    16'h0B0C: data_out = 8'h17;
                    16'h0B0D: data_out = 8'h18;
                    16'h0B0E: data_out = 8'h19;
                    16'h0B0F: data_out = 8'h1A;
                    16'h0B10: data_out = 8'h1B;
                    16'h0B11: data_out = 8'h1C;
                    16'h0B12: data_out = 8'h1D;
                    16'h0B13: data_out = 8'h1E;
                    16'h0B14: data_out = 8'h1F;
                    16'h0B15: data_out = 8'h20;
                    16'h0B16: data_out = 8'h21;
                    16'h0B17: data_out = 8'h22;
                    16'h0B18: data_out = 8'h23;
                    16'h0B19: data_out = 8'h24;
                    16'h0B1A: data_out = 8'h25;
                    16'h0B1B: data_out = 8'h26;
                    16'h0B1C: data_out = 8'h27;
                    16'h0B1D: data_out = 8'h28;
                    16'h0B1E: data_out = 8'h29;
                    16'h0B1F: data_out = 8'h2A;
                    16'h0B20: data_out = 8'h2B;
                    16'h0B21: data_out = 8'h2C;
                    16'h0B22: data_out = 8'h2D;
                    16'h0B23: data_out = 8'h2E;
                    16'h0B24: data_out = 8'h2F;
                    16'h0B25: data_out = 8'h30;
                    16'h0B26: data_out = 8'h31;
                    16'h0B27: data_out = 8'h32;
                    16'h0B28: data_out = 8'h33;
                    16'h0B29: data_out = 8'h34;
                    16'h0B2A: data_out = 8'h35;
                    16'h0B2B: data_out = 8'h36;
                    16'h0B2C: data_out = 8'h37;
                    16'h0B2D: data_out = 8'h38;
                    16'h0B2E: data_out = 8'h39;
                    16'h0B2F: data_out = 8'h3A;
                    16'h0B30: data_out = 8'h3B;
                    16'h0B31: data_out = 8'h3C;
                    16'h0B32: data_out = 8'h3D;
                    16'h0B33: data_out = 8'h3E;
                    16'h0B34: data_out = 8'h3F;
                    16'h0B35: data_out = 8'h40;
                    16'h0B36: data_out = 8'h41;
                    16'h0B37: data_out = 8'h42;
                    16'h0B38: data_out = 8'h43;
                    16'h0B39: data_out = 8'h44;
                    16'h0B3A: data_out = 8'h45;
                    16'h0B3B: data_out = 8'h46;
                    16'h0B3C: data_out = 8'h47;
                    16'h0B3D: data_out = 8'h48;
                    16'h0B3E: data_out = 8'h49;
                    16'h0B3F: data_out = 8'h4A;
                    16'h0B40: data_out = 8'h4B;
                    16'h0B41: data_out = 8'h4C;
                    16'h0B42: data_out = 8'h4D;
                    16'h0B43: data_out = 8'h4E;
                    16'h0B44: data_out = 8'h4F;
                    16'h0B45: data_out = 8'h50;
                    16'h0B46: data_out = 8'h51;
                    16'h0B47: data_out = 8'h52;
                    16'h0B48: data_out = 8'h53;
                    16'h0B49: data_out = 8'h54;
                    16'h0B4A: data_out = 8'h55;
                    16'h0B4B: data_out = 8'h56;
                    16'h0B4C: data_out = 8'h57;
                    16'h0B4D: data_out = 8'h58;
                    16'h0B4E: data_out = 8'h59;
                    16'h0B4F: data_out = 8'h5A;
                    16'h0B50: data_out = 8'h5B;
                    16'h0B51: data_out = 8'h5C;
                    16'h0B52: data_out = 8'h5D;
                    16'h0B53: data_out = 8'h5E;
                    16'h0B54: data_out = 8'h5F;
                    16'h0B55: data_out = 8'h60;
                    16'h0B56: data_out = 8'h61;
                    16'h0B57: data_out = 8'h62;
                    16'h0B58: data_out = 8'h63;
                    16'h0B59: data_out = 8'h64;
                    16'h0B5A: data_out = 8'h65;
                    16'h0B5B: data_out = 8'h66;
                    16'h0B5C: data_out = 8'h67;
                    16'h0B5D: data_out = 8'h68;
                    16'h0B5E: data_out = 8'h69;
                    16'h0B5F: data_out = 8'h6A;
                    16'h0B60: data_out = 8'h6B;
                    16'h0B61: data_out = 8'h6C;
                    16'h0B62: data_out = 8'h6D;
                    16'h0B63: data_out = 8'h6E;
                    16'h0B64: data_out = 8'h6F;
                    16'h0B65: data_out = 8'h70;
                    16'h0B66: data_out = 8'h71;
                    16'h0B67: data_out = 8'h72;
                    16'h0B68: data_out = 8'h73;
                    16'h0B69: data_out = 8'h74;
                    16'h0B6A: data_out = 8'h75;
                    16'h0B6B: data_out = 8'h76;
                    16'h0B6C: data_out = 8'h77;
                    16'h0B6D: data_out = 8'h78;
                    16'h0B6E: data_out = 8'h79;
                    16'h0B6F: data_out = 8'h7A;
                    16'h0B70: data_out = 8'h7B;
                    16'h0B71: data_out = 8'h7C;
                    16'h0B72: data_out = 8'h7D;
                    16'h0B73: data_out = 8'h7E;
                    16'h0B74: data_out = 8'h7F;
                    16'h0B75: data_out = 8'h80;
                    16'h0B76: data_out = 8'h81;
                    16'h0B77: data_out = 8'h82;
                    16'h0B78: data_out = 8'h83;
                    16'h0B79: data_out = 8'h84;
                    16'h0B7A: data_out = 8'h85;
                    16'h0B7B: data_out = 8'h86;
                    16'h0B7C: data_out = 8'h87;
                    16'h0B7D: data_out = 8'h88;
                    16'h0B7E: data_out = 8'h89;
                    16'h0B7F: data_out = 8'h8A;
                    16'h0B80: data_out = 8'hB;
                    16'h0B81: data_out = 8'hA;
                    16'h0B82: data_out = 8'h9;
                    16'h0B83: data_out = 8'h8;
                    16'h0B84: data_out = 8'h7;
                    16'h0B85: data_out = 8'h6;
                    16'h0B86: data_out = 8'h5;
                    16'h0B87: data_out = 8'h4;
                    16'h0B88: data_out = 8'h3;
                    16'h0B89: data_out = 8'h2;
                    16'h0B8A: data_out = 8'h1;
                    16'h0B8B: data_out = 8'h0;
                    16'h0B8C: data_out = 8'h81;
                    16'h0B8D: data_out = 8'h82;
                    16'h0B8E: data_out = 8'h83;
                    16'h0B8F: data_out = 8'h84;
                    16'h0B90: data_out = 8'h85;
                    16'h0B91: data_out = 8'h86;
                    16'h0B92: data_out = 8'h87;
                    16'h0B93: data_out = 8'h88;
                    16'h0B94: data_out = 8'h89;
                    16'h0B95: data_out = 8'h8A;
                    16'h0B96: data_out = 8'h8B;
                    16'h0B97: data_out = 8'h8C;
                    16'h0B98: data_out = 8'h8D;
                    16'h0B99: data_out = 8'h8E;
                    16'h0B9A: data_out = 8'h8F;
                    16'h0B9B: data_out = 8'h90;
                    16'h0B9C: data_out = 8'h91;
                    16'h0B9D: data_out = 8'h92;
                    16'h0B9E: data_out = 8'h93;
                    16'h0B9F: data_out = 8'h94;
                    16'h0BA0: data_out = 8'h95;
                    16'h0BA1: data_out = 8'h96;
                    16'h0BA2: data_out = 8'h97;
                    16'h0BA3: data_out = 8'h98;
                    16'h0BA4: data_out = 8'h99;
                    16'h0BA5: data_out = 8'h9A;
                    16'h0BA6: data_out = 8'h9B;
                    16'h0BA7: data_out = 8'h9C;
                    16'h0BA8: data_out = 8'h9D;
                    16'h0BA9: data_out = 8'h9E;
                    16'h0BAA: data_out = 8'h9F;
                    16'h0BAB: data_out = 8'hA0;
                    16'h0BAC: data_out = 8'hA1;
                    16'h0BAD: data_out = 8'hA2;
                    16'h0BAE: data_out = 8'hA3;
                    16'h0BAF: data_out = 8'hA4;
                    16'h0BB0: data_out = 8'hA5;
                    16'h0BB1: data_out = 8'hA6;
                    16'h0BB2: data_out = 8'hA7;
                    16'h0BB3: data_out = 8'hA8;
                    16'h0BB4: data_out = 8'hA9;
                    16'h0BB5: data_out = 8'hAA;
                    16'h0BB6: data_out = 8'hAB;
                    16'h0BB7: data_out = 8'hAC;
                    16'h0BB8: data_out = 8'hAD;
                    16'h0BB9: data_out = 8'hAE;
                    16'h0BBA: data_out = 8'hAF;
                    16'h0BBB: data_out = 8'hB0;
                    16'h0BBC: data_out = 8'hB1;
                    16'h0BBD: data_out = 8'hB2;
                    16'h0BBE: data_out = 8'hB3;
                    16'h0BBF: data_out = 8'hB4;
                    16'h0BC0: data_out = 8'hB5;
                    16'h0BC1: data_out = 8'hB6;
                    16'h0BC2: data_out = 8'hB7;
                    16'h0BC3: data_out = 8'hB8;
                    16'h0BC4: data_out = 8'hB9;
                    16'h0BC5: data_out = 8'hBA;
                    16'h0BC6: data_out = 8'hBB;
                    16'h0BC7: data_out = 8'hBC;
                    16'h0BC8: data_out = 8'hBD;
                    16'h0BC9: data_out = 8'hBE;
                    16'h0BCA: data_out = 8'hBF;
                    16'h0BCB: data_out = 8'hC0;
                    16'h0BCC: data_out = 8'hC1;
                    16'h0BCD: data_out = 8'hC2;
                    16'h0BCE: data_out = 8'hC3;
                    16'h0BCF: data_out = 8'hC4;
                    16'h0BD0: data_out = 8'hC5;
                    16'h0BD1: data_out = 8'hC6;
                    16'h0BD2: data_out = 8'hC7;
                    16'h0BD3: data_out = 8'hC8;
                    16'h0BD4: data_out = 8'hC9;
                    16'h0BD5: data_out = 8'hCA;
                    16'h0BD6: data_out = 8'hCB;
                    16'h0BD7: data_out = 8'hCC;
                    16'h0BD8: data_out = 8'hCD;
                    16'h0BD9: data_out = 8'hCE;
                    16'h0BDA: data_out = 8'hCF;
                    16'h0BDB: data_out = 8'hD0;
                    16'h0BDC: data_out = 8'hD1;
                    16'h0BDD: data_out = 8'hD2;
                    16'h0BDE: data_out = 8'hD3;
                    16'h0BDF: data_out = 8'hD4;
                    16'h0BE0: data_out = 8'hD5;
                    16'h0BE1: data_out = 8'hD6;
                    16'h0BE2: data_out = 8'hD7;
                    16'h0BE3: data_out = 8'hD8;
                    16'h0BE4: data_out = 8'hD9;
                    16'h0BE5: data_out = 8'hDA;
                    16'h0BE6: data_out = 8'hDB;
                    16'h0BE7: data_out = 8'hDC;
                    16'h0BE8: data_out = 8'hDD;
                    16'h0BE9: data_out = 8'hDE;
                    16'h0BEA: data_out = 8'hDF;
                    16'h0BEB: data_out = 8'hE0;
                    16'h0BEC: data_out = 8'hE1;
                    16'h0BED: data_out = 8'hE2;
                    16'h0BEE: data_out = 8'hE3;
                    16'h0BEF: data_out = 8'hE4;
                    16'h0BF0: data_out = 8'hE5;
                    16'h0BF1: data_out = 8'hE6;
                    16'h0BF2: data_out = 8'hE7;
                    16'h0BF3: data_out = 8'hE8;
                    16'h0BF4: data_out = 8'hE9;
                    16'h0BF5: data_out = 8'hEA;
                    16'h0BF6: data_out = 8'hEB;
                    16'h0BF7: data_out = 8'hEC;
                    16'h0BF8: data_out = 8'hED;
                    16'h0BF9: data_out = 8'hEE;
                    16'h0BFA: data_out = 8'hEF;
                    16'h0BFB: data_out = 8'hF0;
                    16'h0BFC: data_out = 8'hF1;
                    16'h0BFD: data_out = 8'hF2;
                    16'h0BFE: data_out = 8'hF3;
                    16'h0BFF: data_out = 8'hF4;
                    16'h0C00: data_out = 8'hC;
                    16'h0C01: data_out = 8'hD;
                    16'h0C02: data_out = 8'hE;
                    16'h0C03: data_out = 8'hF;
                    16'h0C04: data_out = 8'h10;
                    16'h0C05: data_out = 8'h11;
                    16'h0C06: data_out = 8'h12;
                    16'h0C07: data_out = 8'h13;
                    16'h0C08: data_out = 8'h14;
                    16'h0C09: data_out = 8'h15;
                    16'h0C0A: data_out = 8'h16;
                    16'h0C0B: data_out = 8'h17;
                    16'h0C0C: data_out = 8'h18;
                    16'h0C0D: data_out = 8'h19;
                    16'h0C0E: data_out = 8'h1A;
                    16'h0C0F: data_out = 8'h1B;
                    16'h0C10: data_out = 8'h1C;
                    16'h0C11: data_out = 8'h1D;
                    16'h0C12: data_out = 8'h1E;
                    16'h0C13: data_out = 8'h1F;
                    16'h0C14: data_out = 8'h20;
                    16'h0C15: data_out = 8'h21;
                    16'h0C16: data_out = 8'h22;
                    16'h0C17: data_out = 8'h23;
                    16'h0C18: data_out = 8'h24;
                    16'h0C19: data_out = 8'h25;
                    16'h0C1A: data_out = 8'h26;
                    16'h0C1B: data_out = 8'h27;
                    16'h0C1C: data_out = 8'h28;
                    16'h0C1D: data_out = 8'h29;
                    16'h0C1E: data_out = 8'h2A;
                    16'h0C1F: data_out = 8'h2B;
                    16'h0C20: data_out = 8'h2C;
                    16'h0C21: data_out = 8'h2D;
                    16'h0C22: data_out = 8'h2E;
                    16'h0C23: data_out = 8'h2F;
                    16'h0C24: data_out = 8'h30;
                    16'h0C25: data_out = 8'h31;
                    16'h0C26: data_out = 8'h32;
                    16'h0C27: data_out = 8'h33;
                    16'h0C28: data_out = 8'h34;
                    16'h0C29: data_out = 8'h35;
                    16'h0C2A: data_out = 8'h36;
                    16'h0C2B: data_out = 8'h37;
                    16'h0C2C: data_out = 8'h38;
                    16'h0C2D: data_out = 8'h39;
                    16'h0C2E: data_out = 8'h3A;
                    16'h0C2F: data_out = 8'h3B;
                    16'h0C30: data_out = 8'h3C;
                    16'h0C31: data_out = 8'h3D;
                    16'h0C32: data_out = 8'h3E;
                    16'h0C33: data_out = 8'h3F;
                    16'h0C34: data_out = 8'h40;
                    16'h0C35: data_out = 8'h41;
                    16'h0C36: data_out = 8'h42;
                    16'h0C37: data_out = 8'h43;
                    16'h0C38: data_out = 8'h44;
                    16'h0C39: data_out = 8'h45;
                    16'h0C3A: data_out = 8'h46;
                    16'h0C3B: data_out = 8'h47;
                    16'h0C3C: data_out = 8'h48;
                    16'h0C3D: data_out = 8'h49;
                    16'h0C3E: data_out = 8'h4A;
                    16'h0C3F: data_out = 8'h4B;
                    16'h0C40: data_out = 8'h4C;
                    16'h0C41: data_out = 8'h4D;
                    16'h0C42: data_out = 8'h4E;
                    16'h0C43: data_out = 8'h4F;
                    16'h0C44: data_out = 8'h50;
                    16'h0C45: data_out = 8'h51;
                    16'h0C46: data_out = 8'h52;
                    16'h0C47: data_out = 8'h53;
                    16'h0C48: data_out = 8'h54;
                    16'h0C49: data_out = 8'h55;
                    16'h0C4A: data_out = 8'h56;
                    16'h0C4B: data_out = 8'h57;
                    16'h0C4C: data_out = 8'h58;
                    16'h0C4D: data_out = 8'h59;
                    16'h0C4E: data_out = 8'h5A;
                    16'h0C4F: data_out = 8'h5B;
                    16'h0C50: data_out = 8'h5C;
                    16'h0C51: data_out = 8'h5D;
                    16'h0C52: data_out = 8'h5E;
                    16'h0C53: data_out = 8'h5F;
                    16'h0C54: data_out = 8'h60;
                    16'h0C55: data_out = 8'h61;
                    16'h0C56: data_out = 8'h62;
                    16'h0C57: data_out = 8'h63;
                    16'h0C58: data_out = 8'h64;
                    16'h0C59: data_out = 8'h65;
                    16'h0C5A: data_out = 8'h66;
                    16'h0C5B: data_out = 8'h67;
                    16'h0C5C: data_out = 8'h68;
                    16'h0C5D: data_out = 8'h69;
                    16'h0C5E: data_out = 8'h6A;
                    16'h0C5F: data_out = 8'h6B;
                    16'h0C60: data_out = 8'h6C;
                    16'h0C61: data_out = 8'h6D;
                    16'h0C62: data_out = 8'h6E;
                    16'h0C63: data_out = 8'h6F;
                    16'h0C64: data_out = 8'h70;
                    16'h0C65: data_out = 8'h71;
                    16'h0C66: data_out = 8'h72;
                    16'h0C67: data_out = 8'h73;
                    16'h0C68: data_out = 8'h74;
                    16'h0C69: data_out = 8'h75;
                    16'h0C6A: data_out = 8'h76;
                    16'h0C6B: data_out = 8'h77;
                    16'h0C6C: data_out = 8'h78;
                    16'h0C6D: data_out = 8'h79;
                    16'h0C6E: data_out = 8'h7A;
                    16'h0C6F: data_out = 8'h7B;
                    16'h0C70: data_out = 8'h7C;
                    16'h0C71: data_out = 8'h7D;
                    16'h0C72: data_out = 8'h7E;
                    16'h0C73: data_out = 8'h7F;
                    16'h0C74: data_out = 8'h80;
                    16'h0C75: data_out = 8'h81;
                    16'h0C76: data_out = 8'h82;
                    16'h0C77: data_out = 8'h83;
                    16'h0C78: data_out = 8'h84;
                    16'h0C79: data_out = 8'h85;
                    16'h0C7A: data_out = 8'h86;
                    16'h0C7B: data_out = 8'h87;
                    16'h0C7C: data_out = 8'h88;
                    16'h0C7D: data_out = 8'h89;
                    16'h0C7E: data_out = 8'h8A;
                    16'h0C7F: data_out = 8'h8B;
                    16'h0C80: data_out = 8'hC;
                    16'h0C81: data_out = 8'hB;
                    16'h0C82: data_out = 8'hA;
                    16'h0C83: data_out = 8'h9;
                    16'h0C84: data_out = 8'h8;
                    16'h0C85: data_out = 8'h7;
                    16'h0C86: data_out = 8'h6;
                    16'h0C87: data_out = 8'h5;
                    16'h0C88: data_out = 8'h4;
                    16'h0C89: data_out = 8'h3;
                    16'h0C8A: data_out = 8'h2;
                    16'h0C8B: data_out = 8'h1;
                    16'h0C8C: data_out = 8'h0;
                    16'h0C8D: data_out = 8'h81;
                    16'h0C8E: data_out = 8'h82;
                    16'h0C8F: data_out = 8'h83;
                    16'h0C90: data_out = 8'h84;
                    16'h0C91: data_out = 8'h85;
                    16'h0C92: data_out = 8'h86;
                    16'h0C93: data_out = 8'h87;
                    16'h0C94: data_out = 8'h88;
                    16'h0C95: data_out = 8'h89;
                    16'h0C96: data_out = 8'h8A;
                    16'h0C97: data_out = 8'h8B;
                    16'h0C98: data_out = 8'h8C;
                    16'h0C99: data_out = 8'h8D;
                    16'h0C9A: data_out = 8'h8E;
                    16'h0C9B: data_out = 8'h8F;
                    16'h0C9C: data_out = 8'h90;
                    16'h0C9D: data_out = 8'h91;
                    16'h0C9E: data_out = 8'h92;
                    16'h0C9F: data_out = 8'h93;
                    16'h0CA0: data_out = 8'h94;
                    16'h0CA1: data_out = 8'h95;
                    16'h0CA2: data_out = 8'h96;
                    16'h0CA3: data_out = 8'h97;
                    16'h0CA4: data_out = 8'h98;
                    16'h0CA5: data_out = 8'h99;
                    16'h0CA6: data_out = 8'h9A;
                    16'h0CA7: data_out = 8'h9B;
                    16'h0CA8: data_out = 8'h9C;
                    16'h0CA9: data_out = 8'h9D;
                    16'h0CAA: data_out = 8'h9E;
                    16'h0CAB: data_out = 8'h9F;
                    16'h0CAC: data_out = 8'hA0;
                    16'h0CAD: data_out = 8'hA1;
                    16'h0CAE: data_out = 8'hA2;
                    16'h0CAF: data_out = 8'hA3;
                    16'h0CB0: data_out = 8'hA4;
                    16'h0CB1: data_out = 8'hA5;
                    16'h0CB2: data_out = 8'hA6;
                    16'h0CB3: data_out = 8'hA7;
                    16'h0CB4: data_out = 8'hA8;
                    16'h0CB5: data_out = 8'hA9;
                    16'h0CB6: data_out = 8'hAA;
                    16'h0CB7: data_out = 8'hAB;
                    16'h0CB8: data_out = 8'hAC;
                    16'h0CB9: data_out = 8'hAD;
                    16'h0CBA: data_out = 8'hAE;
                    16'h0CBB: data_out = 8'hAF;
                    16'h0CBC: data_out = 8'hB0;
                    16'h0CBD: data_out = 8'hB1;
                    16'h0CBE: data_out = 8'hB2;
                    16'h0CBF: data_out = 8'hB3;
                    16'h0CC0: data_out = 8'hB4;
                    16'h0CC1: data_out = 8'hB5;
                    16'h0CC2: data_out = 8'hB6;
                    16'h0CC3: data_out = 8'hB7;
                    16'h0CC4: data_out = 8'hB8;
                    16'h0CC5: data_out = 8'hB9;
                    16'h0CC6: data_out = 8'hBA;
                    16'h0CC7: data_out = 8'hBB;
                    16'h0CC8: data_out = 8'hBC;
                    16'h0CC9: data_out = 8'hBD;
                    16'h0CCA: data_out = 8'hBE;
                    16'h0CCB: data_out = 8'hBF;
                    16'h0CCC: data_out = 8'hC0;
                    16'h0CCD: data_out = 8'hC1;
                    16'h0CCE: data_out = 8'hC2;
                    16'h0CCF: data_out = 8'hC3;
                    16'h0CD0: data_out = 8'hC4;
                    16'h0CD1: data_out = 8'hC5;
                    16'h0CD2: data_out = 8'hC6;
                    16'h0CD3: data_out = 8'hC7;
                    16'h0CD4: data_out = 8'hC8;
                    16'h0CD5: data_out = 8'hC9;
                    16'h0CD6: data_out = 8'hCA;
                    16'h0CD7: data_out = 8'hCB;
                    16'h0CD8: data_out = 8'hCC;
                    16'h0CD9: data_out = 8'hCD;
                    16'h0CDA: data_out = 8'hCE;
                    16'h0CDB: data_out = 8'hCF;
                    16'h0CDC: data_out = 8'hD0;
                    16'h0CDD: data_out = 8'hD1;
                    16'h0CDE: data_out = 8'hD2;
                    16'h0CDF: data_out = 8'hD3;
                    16'h0CE0: data_out = 8'hD4;
                    16'h0CE1: data_out = 8'hD5;
                    16'h0CE2: data_out = 8'hD6;
                    16'h0CE3: data_out = 8'hD7;
                    16'h0CE4: data_out = 8'hD8;
                    16'h0CE5: data_out = 8'hD9;
                    16'h0CE6: data_out = 8'hDA;
                    16'h0CE7: data_out = 8'hDB;
                    16'h0CE8: data_out = 8'hDC;
                    16'h0CE9: data_out = 8'hDD;
                    16'h0CEA: data_out = 8'hDE;
                    16'h0CEB: data_out = 8'hDF;
                    16'h0CEC: data_out = 8'hE0;
                    16'h0CED: data_out = 8'hE1;
                    16'h0CEE: data_out = 8'hE2;
                    16'h0CEF: data_out = 8'hE3;
                    16'h0CF0: data_out = 8'hE4;
                    16'h0CF1: data_out = 8'hE5;
                    16'h0CF2: data_out = 8'hE6;
                    16'h0CF3: data_out = 8'hE7;
                    16'h0CF4: data_out = 8'hE8;
                    16'h0CF5: data_out = 8'hE9;
                    16'h0CF6: data_out = 8'hEA;
                    16'h0CF7: data_out = 8'hEB;
                    16'h0CF8: data_out = 8'hEC;
                    16'h0CF9: data_out = 8'hED;
                    16'h0CFA: data_out = 8'hEE;
                    16'h0CFB: data_out = 8'hEF;
                    16'h0CFC: data_out = 8'hF0;
                    16'h0CFD: data_out = 8'hF1;
                    16'h0CFE: data_out = 8'hF2;
                    16'h0CFF: data_out = 8'hF3;
                    16'h0D00: data_out = 8'hD;
                    16'h0D01: data_out = 8'hE;
                    16'h0D02: data_out = 8'hF;
                    16'h0D03: data_out = 8'h10;
                    16'h0D04: data_out = 8'h11;
                    16'h0D05: data_out = 8'h12;
                    16'h0D06: data_out = 8'h13;
                    16'h0D07: data_out = 8'h14;
                    16'h0D08: data_out = 8'h15;
                    16'h0D09: data_out = 8'h16;
                    16'h0D0A: data_out = 8'h17;
                    16'h0D0B: data_out = 8'h18;
                    16'h0D0C: data_out = 8'h19;
                    16'h0D0D: data_out = 8'h1A;
                    16'h0D0E: data_out = 8'h1B;
                    16'h0D0F: data_out = 8'h1C;
                    16'h0D10: data_out = 8'h1D;
                    16'h0D11: data_out = 8'h1E;
                    16'h0D12: data_out = 8'h1F;
                    16'h0D13: data_out = 8'h20;
                    16'h0D14: data_out = 8'h21;
                    16'h0D15: data_out = 8'h22;
                    16'h0D16: data_out = 8'h23;
                    16'h0D17: data_out = 8'h24;
                    16'h0D18: data_out = 8'h25;
                    16'h0D19: data_out = 8'h26;
                    16'h0D1A: data_out = 8'h27;
                    16'h0D1B: data_out = 8'h28;
                    16'h0D1C: data_out = 8'h29;
                    16'h0D1D: data_out = 8'h2A;
                    16'h0D1E: data_out = 8'h2B;
                    16'h0D1F: data_out = 8'h2C;
                    16'h0D20: data_out = 8'h2D;
                    16'h0D21: data_out = 8'h2E;
                    16'h0D22: data_out = 8'h2F;
                    16'h0D23: data_out = 8'h30;
                    16'h0D24: data_out = 8'h31;
                    16'h0D25: data_out = 8'h32;
                    16'h0D26: data_out = 8'h33;
                    16'h0D27: data_out = 8'h34;
                    16'h0D28: data_out = 8'h35;
                    16'h0D29: data_out = 8'h36;
                    16'h0D2A: data_out = 8'h37;
                    16'h0D2B: data_out = 8'h38;
                    16'h0D2C: data_out = 8'h39;
                    16'h0D2D: data_out = 8'h3A;
                    16'h0D2E: data_out = 8'h3B;
                    16'h0D2F: data_out = 8'h3C;
                    16'h0D30: data_out = 8'h3D;
                    16'h0D31: data_out = 8'h3E;
                    16'h0D32: data_out = 8'h3F;
                    16'h0D33: data_out = 8'h40;
                    16'h0D34: data_out = 8'h41;
                    16'h0D35: data_out = 8'h42;
                    16'h0D36: data_out = 8'h43;
                    16'h0D37: data_out = 8'h44;
                    16'h0D38: data_out = 8'h45;
                    16'h0D39: data_out = 8'h46;
                    16'h0D3A: data_out = 8'h47;
                    16'h0D3B: data_out = 8'h48;
                    16'h0D3C: data_out = 8'h49;
                    16'h0D3D: data_out = 8'h4A;
                    16'h0D3E: data_out = 8'h4B;
                    16'h0D3F: data_out = 8'h4C;
                    16'h0D40: data_out = 8'h4D;
                    16'h0D41: data_out = 8'h4E;
                    16'h0D42: data_out = 8'h4F;
                    16'h0D43: data_out = 8'h50;
                    16'h0D44: data_out = 8'h51;
                    16'h0D45: data_out = 8'h52;
                    16'h0D46: data_out = 8'h53;
                    16'h0D47: data_out = 8'h54;
                    16'h0D48: data_out = 8'h55;
                    16'h0D49: data_out = 8'h56;
                    16'h0D4A: data_out = 8'h57;
                    16'h0D4B: data_out = 8'h58;
                    16'h0D4C: data_out = 8'h59;
                    16'h0D4D: data_out = 8'h5A;
                    16'h0D4E: data_out = 8'h5B;
                    16'h0D4F: data_out = 8'h5C;
                    16'h0D50: data_out = 8'h5D;
                    16'h0D51: data_out = 8'h5E;
                    16'h0D52: data_out = 8'h5F;
                    16'h0D53: data_out = 8'h60;
                    16'h0D54: data_out = 8'h61;
                    16'h0D55: data_out = 8'h62;
                    16'h0D56: data_out = 8'h63;
                    16'h0D57: data_out = 8'h64;
                    16'h0D58: data_out = 8'h65;
                    16'h0D59: data_out = 8'h66;
                    16'h0D5A: data_out = 8'h67;
                    16'h0D5B: data_out = 8'h68;
                    16'h0D5C: data_out = 8'h69;
                    16'h0D5D: data_out = 8'h6A;
                    16'h0D5E: data_out = 8'h6B;
                    16'h0D5F: data_out = 8'h6C;
                    16'h0D60: data_out = 8'h6D;
                    16'h0D61: data_out = 8'h6E;
                    16'h0D62: data_out = 8'h6F;
                    16'h0D63: data_out = 8'h70;
                    16'h0D64: data_out = 8'h71;
                    16'h0D65: data_out = 8'h72;
                    16'h0D66: data_out = 8'h73;
                    16'h0D67: data_out = 8'h74;
                    16'h0D68: data_out = 8'h75;
                    16'h0D69: data_out = 8'h76;
                    16'h0D6A: data_out = 8'h77;
                    16'h0D6B: data_out = 8'h78;
                    16'h0D6C: data_out = 8'h79;
                    16'h0D6D: data_out = 8'h7A;
                    16'h0D6E: data_out = 8'h7B;
                    16'h0D6F: data_out = 8'h7C;
                    16'h0D70: data_out = 8'h7D;
                    16'h0D71: data_out = 8'h7E;
                    16'h0D72: data_out = 8'h7F;
                    16'h0D73: data_out = 8'h80;
                    16'h0D74: data_out = 8'h81;
                    16'h0D75: data_out = 8'h82;
                    16'h0D76: data_out = 8'h83;
                    16'h0D77: data_out = 8'h84;
                    16'h0D78: data_out = 8'h85;
                    16'h0D79: data_out = 8'h86;
                    16'h0D7A: data_out = 8'h87;
                    16'h0D7B: data_out = 8'h88;
                    16'h0D7C: data_out = 8'h89;
                    16'h0D7D: data_out = 8'h8A;
                    16'h0D7E: data_out = 8'h8B;
                    16'h0D7F: data_out = 8'h8C;
                    16'h0D80: data_out = 8'hD;
                    16'h0D81: data_out = 8'hC;
                    16'h0D82: data_out = 8'hB;
                    16'h0D83: data_out = 8'hA;
                    16'h0D84: data_out = 8'h9;
                    16'h0D85: data_out = 8'h8;
                    16'h0D86: data_out = 8'h7;
                    16'h0D87: data_out = 8'h6;
                    16'h0D88: data_out = 8'h5;
                    16'h0D89: data_out = 8'h4;
                    16'h0D8A: data_out = 8'h3;
                    16'h0D8B: data_out = 8'h2;
                    16'h0D8C: data_out = 8'h1;
                    16'h0D8D: data_out = 8'h0;
                    16'h0D8E: data_out = 8'h81;
                    16'h0D8F: data_out = 8'h82;
                    16'h0D90: data_out = 8'h83;
                    16'h0D91: data_out = 8'h84;
                    16'h0D92: data_out = 8'h85;
                    16'h0D93: data_out = 8'h86;
                    16'h0D94: data_out = 8'h87;
                    16'h0D95: data_out = 8'h88;
                    16'h0D96: data_out = 8'h89;
                    16'h0D97: data_out = 8'h8A;
                    16'h0D98: data_out = 8'h8B;
                    16'h0D99: data_out = 8'h8C;
                    16'h0D9A: data_out = 8'h8D;
                    16'h0D9B: data_out = 8'h8E;
                    16'h0D9C: data_out = 8'h8F;
                    16'h0D9D: data_out = 8'h90;
                    16'h0D9E: data_out = 8'h91;
                    16'h0D9F: data_out = 8'h92;
                    16'h0DA0: data_out = 8'h93;
                    16'h0DA1: data_out = 8'h94;
                    16'h0DA2: data_out = 8'h95;
                    16'h0DA3: data_out = 8'h96;
                    16'h0DA4: data_out = 8'h97;
                    16'h0DA5: data_out = 8'h98;
                    16'h0DA6: data_out = 8'h99;
                    16'h0DA7: data_out = 8'h9A;
                    16'h0DA8: data_out = 8'h9B;
                    16'h0DA9: data_out = 8'h9C;
                    16'h0DAA: data_out = 8'h9D;
                    16'h0DAB: data_out = 8'h9E;
                    16'h0DAC: data_out = 8'h9F;
                    16'h0DAD: data_out = 8'hA0;
                    16'h0DAE: data_out = 8'hA1;
                    16'h0DAF: data_out = 8'hA2;
                    16'h0DB0: data_out = 8'hA3;
                    16'h0DB1: data_out = 8'hA4;
                    16'h0DB2: data_out = 8'hA5;
                    16'h0DB3: data_out = 8'hA6;
                    16'h0DB4: data_out = 8'hA7;
                    16'h0DB5: data_out = 8'hA8;
                    16'h0DB6: data_out = 8'hA9;
                    16'h0DB7: data_out = 8'hAA;
                    16'h0DB8: data_out = 8'hAB;
                    16'h0DB9: data_out = 8'hAC;
                    16'h0DBA: data_out = 8'hAD;
                    16'h0DBB: data_out = 8'hAE;
                    16'h0DBC: data_out = 8'hAF;
                    16'h0DBD: data_out = 8'hB0;
                    16'h0DBE: data_out = 8'hB1;
                    16'h0DBF: data_out = 8'hB2;
                    16'h0DC0: data_out = 8'hB3;
                    16'h0DC1: data_out = 8'hB4;
                    16'h0DC2: data_out = 8'hB5;
                    16'h0DC3: data_out = 8'hB6;
                    16'h0DC4: data_out = 8'hB7;
                    16'h0DC5: data_out = 8'hB8;
                    16'h0DC6: data_out = 8'hB9;
                    16'h0DC7: data_out = 8'hBA;
                    16'h0DC8: data_out = 8'hBB;
                    16'h0DC9: data_out = 8'hBC;
                    16'h0DCA: data_out = 8'hBD;
                    16'h0DCB: data_out = 8'hBE;
                    16'h0DCC: data_out = 8'hBF;
                    16'h0DCD: data_out = 8'hC0;
                    16'h0DCE: data_out = 8'hC1;
                    16'h0DCF: data_out = 8'hC2;
                    16'h0DD0: data_out = 8'hC3;
                    16'h0DD1: data_out = 8'hC4;
                    16'h0DD2: data_out = 8'hC5;
                    16'h0DD3: data_out = 8'hC6;
                    16'h0DD4: data_out = 8'hC7;
                    16'h0DD5: data_out = 8'hC8;
                    16'h0DD6: data_out = 8'hC9;
                    16'h0DD7: data_out = 8'hCA;
                    16'h0DD8: data_out = 8'hCB;
                    16'h0DD9: data_out = 8'hCC;
                    16'h0DDA: data_out = 8'hCD;
                    16'h0DDB: data_out = 8'hCE;
                    16'h0DDC: data_out = 8'hCF;
                    16'h0DDD: data_out = 8'hD0;
                    16'h0DDE: data_out = 8'hD1;
                    16'h0DDF: data_out = 8'hD2;
                    16'h0DE0: data_out = 8'hD3;
                    16'h0DE1: data_out = 8'hD4;
                    16'h0DE2: data_out = 8'hD5;
                    16'h0DE3: data_out = 8'hD6;
                    16'h0DE4: data_out = 8'hD7;
                    16'h0DE5: data_out = 8'hD8;
                    16'h0DE6: data_out = 8'hD9;
                    16'h0DE7: data_out = 8'hDA;
                    16'h0DE8: data_out = 8'hDB;
                    16'h0DE9: data_out = 8'hDC;
                    16'h0DEA: data_out = 8'hDD;
                    16'h0DEB: data_out = 8'hDE;
                    16'h0DEC: data_out = 8'hDF;
                    16'h0DED: data_out = 8'hE0;
                    16'h0DEE: data_out = 8'hE1;
                    16'h0DEF: data_out = 8'hE2;
                    16'h0DF0: data_out = 8'hE3;
                    16'h0DF1: data_out = 8'hE4;
                    16'h0DF2: data_out = 8'hE5;
                    16'h0DF3: data_out = 8'hE6;
                    16'h0DF4: data_out = 8'hE7;
                    16'h0DF5: data_out = 8'hE8;
                    16'h0DF6: data_out = 8'hE9;
                    16'h0DF7: data_out = 8'hEA;
                    16'h0DF8: data_out = 8'hEB;
                    16'h0DF9: data_out = 8'hEC;
                    16'h0DFA: data_out = 8'hED;
                    16'h0DFB: data_out = 8'hEE;
                    16'h0DFC: data_out = 8'hEF;
                    16'h0DFD: data_out = 8'hF0;
                    16'h0DFE: data_out = 8'hF1;
                    16'h0DFF: data_out = 8'hF2;
                    16'h0E00: data_out = 8'hE;
                    16'h0E01: data_out = 8'hF;
                    16'h0E02: data_out = 8'h10;
                    16'h0E03: data_out = 8'h11;
                    16'h0E04: data_out = 8'h12;
                    16'h0E05: data_out = 8'h13;
                    16'h0E06: data_out = 8'h14;
                    16'h0E07: data_out = 8'h15;
                    16'h0E08: data_out = 8'h16;
                    16'h0E09: data_out = 8'h17;
                    16'h0E0A: data_out = 8'h18;
                    16'h0E0B: data_out = 8'h19;
                    16'h0E0C: data_out = 8'h1A;
                    16'h0E0D: data_out = 8'h1B;
                    16'h0E0E: data_out = 8'h1C;
                    16'h0E0F: data_out = 8'h1D;
                    16'h0E10: data_out = 8'h1E;
                    16'h0E11: data_out = 8'h1F;
                    16'h0E12: data_out = 8'h20;
                    16'h0E13: data_out = 8'h21;
                    16'h0E14: data_out = 8'h22;
                    16'h0E15: data_out = 8'h23;
                    16'h0E16: data_out = 8'h24;
                    16'h0E17: data_out = 8'h25;
                    16'h0E18: data_out = 8'h26;
                    16'h0E19: data_out = 8'h27;
                    16'h0E1A: data_out = 8'h28;
                    16'h0E1B: data_out = 8'h29;
                    16'h0E1C: data_out = 8'h2A;
                    16'h0E1D: data_out = 8'h2B;
                    16'h0E1E: data_out = 8'h2C;
                    16'h0E1F: data_out = 8'h2D;
                    16'h0E20: data_out = 8'h2E;
                    16'h0E21: data_out = 8'h2F;
                    16'h0E22: data_out = 8'h30;
                    16'h0E23: data_out = 8'h31;
                    16'h0E24: data_out = 8'h32;
                    16'h0E25: data_out = 8'h33;
                    16'h0E26: data_out = 8'h34;
                    16'h0E27: data_out = 8'h35;
                    16'h0E28: data_out = 8'h36;
                    16'h0E29: data_out = 8'h37;
                    16'h0E2A: data_out = 8'h38;
                    16'h0E2B: data_out = 8'h39;
                    16'h0E2C: data_out = 8'h3A;
                    16'h0E2D: data_out = 8'h3B;
                    16'h0E2E: data_out = 8'h3C;
                    16'h0E2F: data_out = 8'h3D;
                    16'h0E30: data_out = 8'h3E;
                    16'h0E31: data_out = 8'h3F;
                    16'h0E32: data_out = 8'h40;
                    16'h0E33: data_out = 8'h41;
                    16'h0E34: data_out = 8'h42;
                    16'h0E35: data_out = 8'h43;
                    16'h0E36: data_out = 8'h44;
                    16'h0E37: data_out = 8'h45;
                    16'h0E38: data_out = 8'h46;
                    16'h0E39: data_out = 8'h47;
                    16'h0E3A: data_out = 8'h48;
                    16'h0E3B: data_out = 8'h49;
                    16'h0E3C: data_out = 8'h4A;
                    16'h0E3D: data_out = 8'h4B;
                    16'h0E3E: data_out = 8'h4C;
                    16'h0E3F: data_out = 8'h4D;
                    16'h0E40: data_out = 8'h4E;
                    16'h0E41: data_out = 8'h4F;
                    16'h0E42: data_out = 8'h50;
                    16'h0E43: data_out = 8'h51;
                    16'h0E44: data_out = 8'h52;
                    16'h0E45: data_out = 8'h53;
                    16'h0E46: data_out = 8'h54;
                    16'h0E47: data_out = 8'h55;
                    16'h0E48: data_out = 8'h56;
                    16'h0E49: data_out = 8'h57;
                    16'h0E4A: data_out = 8'h58;
                    16'h0E4B: data_out = 8'h59;
                    16'h0E4C: data_out = 8'h5A;
                    16'h0E4D: data_out = 8'h5B;
                    16'h0E4E: data_out = 8'h5C;
                    16'h0E4F: data_out = 8'h5D;
                    16'h0E50: data_out = 8'h5E;
                    16'h0E51: data_out = 8'h5F;
                    16'h0E52: data_out = 8'h60;
                    16'h0E53: data_out = 8'h61;
                    16'h0E54: data_out = 8'h62;
                    16'h0E55: data_out = 8'h63;
                    16'h0E56: data_out = 8'h64;
                    16'h0E57: data_out = 8'h65;
                    16'h0E58: data_out = 8'h66;
                    16'h0E59: data_out = 8'h67;
                    16'h0E5A: data_out = 8'h68;
                    16'h0E5B: data_out = 8'h69;
                    16'h0E5C: data_out = 8'h6A;
                    16'h0E5D: data_out = 8'h6B;
                    16'h0E5E: data_out = 8'h6C;
                    16'h0E5F: data_out = 8'h6D;
                    16'h0E60: data_out = 8'h6E;
                    16'h0E61: data_out = 8'h6F;
                    16'h0E62: data_out = 8'h70;
                    16'h0E63: data_out = 8'h71;
                    16'h0E64: data_out = 8'h72;
                    16'h0E65: data_out = 8'h73;
                    16'h0E66: data_out = 8'h74;
                    16'h0E67: data_out = 8'h75;
                    16'h0E68: data_out = 8'h76;
                    16'h0E69: data_out = 8'h77;
                    16'h0E6A: data_out = 8'h78;
                    16'h0E6B: data_out = 8'h79;
                    16'h0E6C: data_out = 8'h7A;
                    16'h0E6D: data_out = 8'h7B;
                    16'h0E6E: data_out = 8'h7C;
                    16'h0E6F: data_out = 8'h7D;
                    16'h0E70: data_out = 8'h7E;
                    16'h0E71: data_out = 8'h7F;
                    16'h0E72: data_out = 8'h80;
                    16'h0E73: data_out = 8'h81;
                    16'h0E74: data_out = 8'h82;
                    16'h0E75: data_out = 8'h83;
                    16'h0E76: data_out = 8'h84;
                    16'h0E77: data_out = 8'h85;
                    16'h0E78: data_out = 8'h86;
                    16'h0E79: data_out = 8'h87;
                    16'h0E7A: data_out = 8'h88;
                    16'h0E7B: data_out = 8'h89;
                    16'h0E7C: data_out = 8'h8A;
                    16'h0E7D: data_out = 8'h8B;
                    16'h0E7E: data_out = 8'h8C;
                    16'h0E7F: data_out = 8'h8D;
                    16'h0E80: data_out = 8'hE;
                    16'h0E81: data_out = 8'hD;
                    16'h0E82: data_out = 8'hC;
                    16'h0E83: data_out = 8'hB;
                    16'h0E84: data_out = 8'hA;
                    16'h0E85: data_out = 8'h9;
                    16'h0E86: data_out = 8'h8;
                    16'h0E87: data_out = 8'h7;
                    16'h0E88: data_out = 8'h6;
                    16'h0E89: data_out = 8'h5;
                    16'h0E8A: data_out = 8'h4;
                    16'h0E8B: data_out = 8'h3;
                    16'h0E8C: data_out = 8'h2;
                    16'h0E8D: data_out = 8'h1;
                    16'h0E8E: data_out = 8'h0;
                    16'h0E8F: data_out = 8'h81;
                    16'h0E90: data_out = 8'h82;
                    16'h0E91: data_out = 8'h83;
                    16'h0E92: data_out = 8'h84;
                    16'h0E93: data_out = 8'h85;
                    16'h0E94: data_out = 8'h86;
                    16'h0E95: data_out = 8'h87;
                    16'h0E96: data_out = 8'h88;
                    16'h0E97: data_out = 8'h89;
                    16'h0E98: data_out = 8'h8A;
                    16'h0E99: data_out = 8'h8B;
                    16'h0E9A: data_out = 8'h8C;
                    16'h0E9B: data_out = 8'h8D;
                    16'h0E9C: data_out = 8'h8E;
                    16'h0E9D: data_out = 8'h8F;
                    16'h0E9E: data_out = 8'h90;
                    16'h0E9F: data_out = 8'h91;
                    16'h0EA0: data_out = 8'h92;
                    16'h0EA1: data_out = 8'h93;
                    16'h0EA2: data_out = 8'h94;
                    16'h0EA3: data_out = 8'h95;
                    16'h0EA4: data_out = 8'h96;
                    16'h0EA5: data_out = 8'h97;
                    16'h0EA6: data_out = 8'h98;
                    16'h0EA7: data_out = 8'h99;
                    16'h0EA8: data_out = 8'h9A;
                    16'h0EA9: data_out = 8'h9B;
                    16'h0EAA: data_out = 8'h9C;
                    16'h0EAB: data_out = 8'h9D;
                    16'h0EAC: data_out = 8'h9E;
                    16'h0EAD: data_out = 8'h9F;
                    16'h0EAE: data_out = 8'hA0;
                    16'h0EAF: data_out = 8'hA1;
                    16'h0EB0: data_out = 8'hA2;
                    16'h0EB1: data_out = 8'hA3;
                    16'h0EB2: data_out = 8'hA4;
                    16'h0EB3: data_out = 8'hA5;
                    16'h0EB4: data_out = 8'hA6;
                    16'h0EB5: data_out = 8'hA7;
                    16'h0EB6: data_out = 8'hA8;
                    16'h0EB7: data_out = 8'hA9;
                    16'h0EB8: data_out = 8'hAA;
                    16'h0EB9: data_out = 8'hAB;
                    16'h0EBA: data_out = 8'hAC;
                    16'h0EBB: data_out = 8'hAD;
                    16'h0EBC: data_out = 8'hAE;
                    16'h0EBD: data_out = 8'hAF;
                    16'h0EBE: data_out = 8'hB0;
                    16'h0EBF: data_out = 8'hB1;
                    16'h0EC0: data_out = 8'hB2;
                    16'h0EC1: data_out = 8'hB3;
                    16'h0EC2: data_out = 8'hB4;
                    16'h0EC3: data_out = 8'hB5;
                    16'h0EC4: data_out = 8'hB6;
                    16'h0EC5: data_out = 8'hB7;
                    16'h0EC6: data_out = 8'hB8;
                    16'h0EC7: data_out = 8'hB9;
                    16'h0EC8: data_out = 8'hBA;
                    16'h0EC9: data_out = 8'hBB;
                    16'h0ECA: data_out = 8'hBC;
                    16'h0ECB: data_out = 8'hBD;
                    16'h0ECC: data_out = 8'hBE;
                    16'h0ECD: data_out = 8'hBF;
                    16'h0ECE: data_out = 8'hC0;
                    16'h0ECF: data_out = 8'hC1;
                    16'h0ED0: data_out = 8'hC2;
                    16'h0ED1: data_out = 8'hC3;
                    16'h0ED2: data_out = 8'hC4;
                    16'h0ED3: data_out = 8'hC5;
                    16'h0ED4: data_out = 8'hC6;
                    16'h0ED5: data_out = 8'hC7;
                    16'h0ED6: data_out = 8'hC8;
                    16'h0ED7: data_out = 8'hC9;
                    16'h0ED8: data_out = 8'hCA;
                    16'h0ED9: data_out = 8'hCB;
                    16'h0EDA: data_out = 8'hCC;
                    16'h0EDB: data_out = 8'hCD;
                    16'h0EDC: data_out = 8'hCE;
                    16'h0EDD: data_out = 8'hCF;
                    16'h0EDE: data_out = 8'hD0;
                    16'h0EDF: data_out = 8'hD1;
                    16'h0EE0: data_out = 8'hD2;
                    16'h0EE1: data_out = 8'hD3;
                    16'h0EE2: data_out = 8'hD4;
                    16'h0EE3: data_out = 8'hD5;
                    16'h0EE4: data_out = 8'hD6;
                    16'h0EE5: data_out = 8'hD7;
                    16'h0EE6: data_out = 8'hD8;
                    16'h0EE7: data_out = 8'hD9;
                    16'h0EE8: data_out = 8'hDA;
                    16'h0EE9: data_out = 8'hDB;
                    16'h0EEA: data_out = 8'hDC;
                    16'h0EEB: data_out = 8'hDD;
                    16'h0EEC: data_out = 8'hDE;
                    16'h0EED: data_out = 8'hDF;
                    16'h0EEE: data_out = 8'hE0;
                    16'h0EEF: data_out = 8'hE1;
                    16'h0EF0: data_out = 8'hE2;
                    16'h0EF1: data_out = 8'hE3;
                    16'h0EF2: data_out = 8'hE4;
                    16'h0EF3: data_out = 8'hE5;
                    16'h0EF4: data_out = 8'hE6;
                    16'h0EF5: data_out = 8'hE7;
                    16'h0EF6: data_out = 8'hE8;
                    16'h0EF7: data_out = 8'hE9;
                    16'h0EF8: data_out = 8'hEA;
                    16'h0EF9: data_out = 8'hEB;
                    16'h0EFA: data_out = 8'hEC;
                    16'h0EFB: data_out = 8'hED;
                    16'h0EFC: data_out = 8'hEE;
                    16'h0EFD: data_out = 8'hEF;
                    16'h0EFE: data_out = 8'hF0;
                    16'h0EFF: data_out = 8'hF1;
                    16'h0F00: data_out = 8'hF;
                    16'h0F01: data_out = 8'h10;
                    16'h0F02: data_out = 8'h11;
                    16'h0F03: data_out = 8'h12;
                    16'h0F04: data_out = 8'h13;
                    16'h0F05: data_out = 8'h14;
                    16'h0F06: data_out = 8'h15;
                    16'h0F07: data_out = 8'h16;
                    16'h0F08: data_out = 8'h17;
                    16'h0F09: data_out = 8'h18;
                    16'h0F0A: data_out = 8'h19;
                    16'h0F0B: data_out = 8'h1A;
                    16'h0F0C: data_out = 8'h1B;
                    16'h0F0D: data_out = 8'h1C;
                    16'h0F0E: data_out = 8'h1D;
                    16'h0F0F: data_out = 8'h1E;
                    16'h0F10: data_out = 8'h1F;
                    16'h0F11: data_out = 8'h20;
                    16'h0F12: data_out = 8'h21;
                    16'h0F13: data_out = 8'h22;
                    16'h0F14: data_out = 8'h23;
                    16'h0F15: data_out = 8'h24;
                    16'h0F16: data_out = 8'h25;
                    16'h0F17: data_out = 8'h26;
                    16'h0F18: data_out = 8'h27;
                    16'h0F19: data_out = 8'h28;
                    16'h0F1A: data_out = 8'h29;
                    16'h0F1B: data_out = 8'h2A;
                    16'h0F1C: data_out = 8'h2B;
                    16'h0F1D: data_out = 8'h2C;
                    16'h0F1E: data_out = 8'h2D;
                    16'h0F1F: data_out = 8'h2E;
                    16'h0F20: data_out = 8'h2F;
                    16'h0F21: data_out = 8'h30;
                    16'h0F22: data_out = 8'h31;
                    16'h0F23: data_out = 8'h32;
                    16'h0F24: data_out = 8'h33;
                    16'h0F25: data_out = 8'h34;
                    16'h0F26: data_out = 8'h35;
                    16'h0F27: data_out = 8'h36;
                    16'h0F28: data_out = 8'h37;
                    16'h0F29: data_out = 8'h38;
                    16'h0F2A: data_out = 8'h39;
                    16'h0F2B: data_out = 8'h3A;
                    16'h0F2C: data_out = 8'h3B;
                    16'h0F2D: data_out = 8'h3C;
                    16'h0F2E: data_out = 8'h3D;
                    16'h0F2F: data_out = 8'h3E;
                    16'h0F30: data_out = 8'h3F;
                    16'h0F31: data_out = 8'h40;
                    16'h0F32: data_out = 8'h41;
                    16'h0F33: data_out = 8'h42;
                    16'h0F34: data_out = 8'h43;
                    16'h0F35: data_out = 8'h44;
                    16'h0F36: data_out = 8'h45;
                    16'h0F37: data_out = 8'h46;
                    16'h0F38: data_out = 8'h47;
                    16'h0F39: data_out = 8'h48;
                    16'h0F3A: data_out = 8'h49;
                    16'h0F3B: data_out = 8'h4A;
                    16'h0F3C: data_out = 8'h4B;
                    16'h0F3D: data_out = 8'h4C;
                    16'h0F3E: data_out = 8'h4D;
                    16'h0F3F: data_out = 8'h4E;
                    16'h0F40: data_out = 8'h4F;
                    16'h0F41: data_out = 8'h50;
                    16'h0F42: data_out = 8'h51;
                    16'h0F43: data_out = 8'h52;
                    16'h0F44: data_out = 8'h53;
                    16'h0F45: data_out = 8'h54;
                    16'h0F46: data_out = 8'h55;
                    16'h0F47: data_out = 8'h56;
                    16'h0F48: data_out = 8'h57;
                    16'h0F49: data_out = 8'h58;
                    16'h0F4A: data_out = 8'h59;
                    16'h0F4B: data_out = 8'h5A;
                    16'h0F4C: data_out = 8'h5B;
                    16'h0F4D: data_out = 8'h5C;
                    16'h0F4E: data_out = 8'h5D;
                    16'h0F4F: data_out = 8'h5E;
                    16'h0F50: data_out = 8'h5F;
                    16'h0F51: data_out = 8'h60;
                    16'h0F52: data_out = 8'h61;
                    16'h0F53: data_out = 8'h62;
                    16'h0F54: data_out = 8'h63;
                    16'h0F55: data_out = 8'h64;
                    16'h0F56: data_out = 8'h65;
                    16'h0F57: data_out = 8'h66;
                    16'h0F58: data_out = 8'h67;
                    16'h0F59: data_out = 8'h68;
                    16'h0F5A: data_out = 8'h69;
                    16'h0F5B: data_out = 8'h6A;
                    16'h0F5C: data_out = 8'h6B;
                    16'h0F5D: data_out = 8'h6C;
                    16'h0F5E: data_out = 8'h6D;
                    16'h0F5F: data_out = 8'h6E;
                    16'h0F60: data_out = 8'h6F;
                    16'h0F61: data_out = 8'h70;
                    16'h0F62: data_out = 8'h71;
                    16'h0F63: data_out = 8'h72;
                    16'h0F64: data_out = 8'h73;
                    16'h0F65: data_out = 8'h74;
                    16'h0F66: data_out = 8'h75;
                    16'h0F67: data_out = 8'h76;
                    16'h0F68: data_out = 8'h77;
                    16'h0F69: data_out = 8'h78;
                    16'h0F6A: data_out = 8'h79;
                    16'h0F6B: data_out = 8'h7A;
                    16'h0F6C: data_out = 8'h7B;
                    16'h0F6D: data_out = 8'h7C;
                    16'h0F6E: data_out = 8'h7D;
                    16'h0F6F: data_out = 8'h7E;
                    16'h0F70: data_out = 8'h7F;
                    16'h0F71: data_out = 8'h80;
                    16'h0F72: data_out = 8'h81;
                    16'h0F73: data_out = 8'h82;
                    16'h0F74: data_out = 8'h83;
                    16'h0F75: data_out = 8'h84;
                    16'h0F76: data_out = 8'h85;
                    16'h0F77: data_out = 8'h86;
                    16'h0F78: data_out = 8'h87;
                    16'h0F79: data_out = 8'h88;
                    16'h0F7A: data_out = 8'h89;
                    16'h0F7B: data_out = 8'h8A;
                    16'h0F7C: data_out = 8'h8B;
                    16'h0F7D: data_out = 8'h8C;
                    16'h0F7E: data_out = 8'h8D;
                    16'h0F7F: data_out = 8'h8E;
                    16'h0F80: data_out = 8'hF;
                    16'h0F81: data_out = 8'hE;
                    16'h0F82: data_out = 8'hD;
                    16'h0F83: data_out = 8'hC;
                    16'h0F84: data_out = 8'hB;
                    16'h0F85: data_out = 8'hA;
                    16'h0F86: data_out = 8'h9;
                    16'h0F87: data_out = 8'h8;
                    16'h0F88: data_out = 8'h7;
                    16'h0F89: data_out = 8'h6;
                    16'h0F8A: data_out = 8'h5;
                    16'h0F8B: data_out = 8'h4;
                    16'h0F8C: data_out = 8'h3;
                    16'h0F8D: data_out = 8'h2;
                    16'h0F8E: data_out = 8'h1;
                    16'h0F8F: data_out = 8'h0;
                    16'h0F90: data_out = 8'h81;
                    16'h0F91: data_out = 8'h82;
                    16'h0F92: data_out = 8'h83;
                    16'h0F93: data_out = 8'h84;
                    16'h0F94: data_out = 8'h85;
                    16'h0F95: data_out = 8'h86;
                    16'h0F96: data_out = 8'h87;
                    16'h0F97: data_out = 8'h88;
                    16'h0F98: data_out = 8'h89;
                    16'h0F99: data_out = 8'h8A;
                    16'h0F9A: data_out = 8'h8B;
                    16'h0F9B: data_out = 8'h8C;
                    16'h0F9C: data_out = 8'h8D;
                    16'h0F9D: data_out = 8'h8E;
                    16'h0F9E: data_out = 8'h8F;
                    16'h0F9F: data_out = 8'h90;
                    16'h0FA0: data_out = 8'h91;
                    16'h0FA1: data_out = 8'h92;
                    16'h0FA2: data_out = 8'h93;
                    16'h0FA3: data_out = 8'h94;
                    16'h0FA4: data_out = 8'h95;
                    16'h0FA5: data_out = 8'h96;
                    16'h0FA6: data_out = 8'h97;
                    16'h0FA7: data_out = 8'h98;
                    16'h0FA8: data_out = 8'h99;
                    16'h0FA9: data_out = 8'h9A;
                    16'h0FAA: data_out = 8'h9B;
                    16'h0FAB: data_out = 8'h9C;
                    16'h0FAC: data_out = 8'h9D;
                    16'h0FAD: data_out = 8'h9E;
                    16'h0FAE: data_out = 8'h9F;
                    16'h0FAF: data_out = 8'hA0;
                    16'h0FB0: data_out = 8'hA1;
                    16'h0FB1: data_out = 8'hA2;
                    16'h0FB2: data_out = 8'hA3;
                    16'h0FB3: data_out = 8'hA4;
                    16'h0FB4: data_out = 8'hA5;
                    16'h0FB5: data_out = 8'hA6;
                    16'h0FB6: data_out = 8'hA7;
                    16'h0FB7: data_out = 8'hA8;
                    16'h0FB8: data_out = 8'hA9;
                    16'h0FB9: data_out = 8'hAA;
                    16'h0FBA: data_out = 8'hAB;
                    16'h0FBB: data_out = 8'hAC;
                    16'h0FBC: data_out = 8'hAD;
                    16'h0FBD: data_out = 8'hAE;
                    16'h0FBE: data_out = 8'hAF;
                    16'h0FBF: data_out = 8'hB0;
                    16'h0FC0: data_out = 8'hB1;
                    16'h0FC1: data_out = 8'hB2;
                    16'h0FC2: data_out = 8'hB3;
                    16'h0FC3: data_out = 8'hB4;
                    16'h0FC4: data_out = 8'hB5;
                    16'h0FC5: data_out = 8'hB6;
                    16'h0FC6: data_out = 8'hB7;
                    16'h0FC7: data_out = 8'hB8;
                    16'h0FC8: data_out = 8'hB9;
                    16'h0FC9: data_out = 8'hBA;
                    16'h0FCA: data_out = 8'hBB;
                    16'h0FCB: data_out = 8'hBC;
                    16'h0FCC: data_out = 8'hBD;
                    16'h0FCD: data_out = 8'hBE;
                    16'h0FCE: data_out = 8'hBF;
                    16'h0FCF: data_out = 8'hC0;
                    16'h0FD0: data_out = 8'hC1;
                    16'h0FD1: data_out = 8'hC2;
                    16'h0FD2: data_out = 8'hC3;
                    16'h0FD3: data_out = 8'hC4;
                    16'h0FD4: data_out = 8'hC5;
                    16'h0FD5: data_out = 8'hC6;
                    16'h0FD6: data_out = 8'hC7;
                    16'h0FD7: data_out = 8'hC8;
                    16'h0FD8: data_out = 8'hC9;
                    16'h0FD9: data_out = 8'hCA;
                    16'h0FDA: data_out = 8'hCB;
                    16'h0FDB: data_out = 8'hCC;
                    16'h0FDC: data_out = 8'hCD;
                    16'h0FDD: data_out = 8'hCE;
                    16'h0FDE: data_out = 8'hCF;
                    16'h0FDF: data_out = 8'hD0;
                    16'h0FE0: data_out = 8'hD1;
                    16'h0FE1: data_out = 8'hD2;
                    16'h0FE2: data_out = 8'hD3;
                    16'h0FE3: data_out = 8'hD4;
                    16'h0FE4: data_out = 8'hD5;
                    16'h0FE5: data_out = 8'hD6;
                    16'h0FE6: data_out = 8'hD7;
                    16'h0FE7: data_out = 8'hD8;
                    16'h0FE8: data_out = 8'hD9;
                    16'h0FE9: data_out = 8'hDA;
                    16'h0FEA: data_out = 8'hDB;
                    16'h0FEB: data_out = 8'hDC;
                    16'h0FEC: data_out = 8'hDD;
                    16'h0FED: data_out = 8'hDE;
                    16'h0FEE: data_out = 8'hDF;
                    16'h0FEF: data_out = 8'hE0;
                    16'h0FF0: data_out = 8'hE1;
                    16'h0FF1: data_out = 8'hE2;
                    16'h0FF2: data_out = 8'hE3;
                    16'h0FF3: data_out = 8'hE4;
                    16'h0FF4: data_out = 8'hE5;
                    16'h0FF5: data_out = 8'hE6;
                    16'h0FF6: data_out = 8'hE7;
                    16'h0FF7: data_out = 8'hE8;
                    16'h0FF8: data_out = 8'hE9;
                    16'h0FF9: data_out = 8'hEA;
                    16'h0FFA: data_out = 8'hEB;
                    16'h0FFB: data_out = 8'hEC;
                    16'h0FFC: data_out = 8'hED;
                    16'h0FFD: data_out = 8'hEE;
                    16'h0FFE: data_out = 8'hEF;
                    16'h0FFF: data_out = 8'hF0;
                    16'h1000: data_out = 8'h10;
                    16'h1001: data_out = 8'h11;
                    16'h1002: data_out = 8'h12;
                    16'h1003: data_out = 8'h13;
                    16'h1004: data_out = 8'h14;
                    16'h1005: data_out = 8'h15;
                    16'h1006: data_out = 8'h16;
                    16'h1007: data_out = 8'h17;
                    16'h1008: data_out = 8'h18;
                    16'h1009: data_out = 8'h19;
                    16'h100A: data_out = 8'h1A;
                    16'h100B: data_out = 8'h1B;
                    16'h100C: data_out = 8'h1C;
                    16'h100D: data_out = 8'h1D;
                    16'h100E: data_out = 8'h1E;
                    16'h100F: data_out = 8'h1F;
                    16'h1010: data_out = 8'h20;
                    16'h1011: data_out = 8'h21;
                    16'h1012: data_out = 8'h22;
                    16'h1013: data_out = 8'h23;
                    16'h1014: data_out = 8'h24;
                    16'h1015: data_out = 8'h25;
                    16'h1016: data_out = 8'h26;
                    16'h1017: data_out = 8'h27;
                    16'h1018: data_out = 8'h28;
                    16'h1019: data_out = 8'h29;
                    16'h101A: data_out = 8'h2A;
                    16'h101B: data_out = 8'h2B;
                    16'h101C: data_out = 8'h2C;
                    16'h101D: data_out = 8'h2D;
                    16'h101E: data_out = 8'h2E;
                    16'h101F: data_out = 8'h2F;
                    16'h1020: data_out = 8'h30;
                    16'h1021: data_out = 8'h31;
                    16'h1022: data_out = 8'h32;
                    16'h1023: data_out = 8'h33;
                    16'h1024: data_out = 8'h34;
                    16'h1025: data_out = 8'h35;
                    16'h1026: data_out = 8'h36;
                    16'h1027: data_out = 8'h37;
                    16'h1028: data_out = 8'h38;
                    16'h1029: data_out = 8'h39;
                    16'h102A: data_out = 8'h3A;
                    16'h102B: data_out = 8'h3B;
                    16'h102C: data_out = 8'h3C;
                    16'h102D: data_out = 8'h3D;
                    16'h102E: data_out = 8'h3E;
                    16'h102F: data_out = 8'h3F;
                    16'h1030: data_out = 8'h40;
                    16'h1031: data_out = 8'h41;
                    16'h1032: data_out = 8'h42;
                    16'h1033: data_out = 8'h43;
                    16'h1034: data_out = 8'h44;
                    16'h1035: data_out = 8'h45;
                    16'h1036: data_out = 8'h46;
                    16'h1037: data_out = 8'h47;
                    16'h1038: data_out = 8'h48;
                    16'h1039: data_out = 8'h49;
                    16'h103A: data_out = 8'h4A;
                    16'h103B: data_out = 8'h4B;
                    16'h103C: data_out = 8'h4C;
                    16'h103D: data_out = 8'h4D;
                    16'h103E: data_out = 8'h4E;
                    16'h103F: data_out = 8'h4F;
                    16'h1040: data_out = 8'h50;
                    16'h1041: data_out = 8'h51;
                    16'h1042: data_out = 8'h52;
                    16'h1043: data_out = 8'h53;
                    16'h1044: data_out = 8'h54;
                    16'h1045: data_out = 8'h55;
                    16'h1046: data_out = 8'h56;
                    16'h1047: data_out = 8'h57;
                    16'h1048: data_out = 8'h58;
                    16'h1049: data_out = 8'h59;
                    16'h104A: data_out = 8'h5A;
                    16'h104B: data_out = 8'h5B;
                    16'h104C: data_out = 8'h5C;
                    16'h104D: data_out = 8'h5D;
                    16'h104E: data_out = 8'h5E;
                    16'h104F: data_out = 8'h5F;
                    16'h1050: data_out = 8'h60;
                    16'h1051: data_out = 8'h61;
                    16'h1052: data_out = 8'h62;
                    16'h1053: data_out = 8'h63;
                    16'h1054: data_out = 8'h64;
                    16'h1055: data_out = 8'h65;
                    16'h1056: data_out = 8'h66;
                    16'h1057: data_out = 8'h67;
                    16'h1058: data_out = 8'h68;
                    16'h1059: data_out = 8'h69;
                    16'h105A: data_out = 8'h6A;
                    16'h105B: data_out = 8'h6B;
                    16'h105C: data_out = 8'h6C;
                    16'h105D: data_out = 8'h6D;
                    16'h105E: data_out = 8'h6E;
                    16'h105F: data_out = 8'h6F;
                    16'h1060: data_out = 8'h70;
                    16'h1061: data_out = 8'h71;
                    16'h1062: data_out = 8'h72;
                    16'h1063: data_out = 8'h73;
                    16'h1064: data_out = 8'h74;
                    16'h1065: data_out = 8'h75;
                    16'h1066: data_out = 8'h76;
                    16'h1067: data_out = 8'h77;
                    16'h1068: data_out = 8'h78;
                    16'h1069: data_out = 8'h79;
                    16'h106A: data_out = 8'h7A;
                    16'h106B: data_out = 8'h7B;
                    16'h106C: data_out = 8'h7C;
                    16'h106D: data_out = 8'h7D;
                    16'h106E: data_out = 8'h7E;
                    16'h106F: data_out = 8'h7F;
                    16'h1070: data_out = 8'h80;
                    16'h1071: data_out = 8'h81;
                    16'h1072: data_out = 8'h82;
                    16'h1073: data_out = 8'h83;
                    16'h1074: data_out = 8'h84;
                    16'h1075: data_out = 8'h85;
                    16'h1076: data_out = 8'h86;
                    16'h1077: data_out = 8'h87;
                    16'h1078: data_out = 8'h88;
                    16'h1079: data_out = 8'h89;
                    16'h107A: data_out = 8'h8A;
                    16'h107B: data_out = 8'h8B;
                    16'h107C: data_out = 8'h8C;
                    16'h107D: data_out = 8'h8D;
                    16'h107E: data_out = 8'h8E;
                    16'h107F: data_out = 8'h8F;
                    16'h1080: data_out = 8'h10;
                    16'h1081: data_out = 8'hF;
                    16'h1082: data_out = 8'hE;
                    16'h1083: data_out = 8'hD;
                    16'h1084: data_out = 8'hC;
                    16'h1085: data_out = 8'hB;
                    16'h1086: data_out = 8'hA;
                    16'h1087: data_out = 8'h9;
                    16'h1088: data_out = 8'h8;
                    16'h1089: data_out = 8'h7;
                    16'h108A: data_out = 8'h6;
                    16'h108B: data_out = 8'h5;
                    16'h108C: data_out = 8'h4;
                    16'h108D: data_out = 8'h3;
                    16'h108E: data_out = 8'h2;
                    16'h108F: data_out = 8'h1;
                    16'h1090: data_out = 8'h0;
                    16'h1091: data_out = 8'h81;
                    16'h1092: data_out = 8'h82;
                    16'h1093: data_out = 8'h83;
                    16'h1094: data_out = 8'h84;
                    16'h1095: data_out = 8'h85;
                    16'h1096: data_out = 8'h86;
                    16'h1097: data_out = 8'h87;
                    16'h1098: data_out = 8'h88;
                    16'h1099: data_out = 8'h89;
                    16'h109A: data_out = 8'h8A;
                    16'h109B: data_out = 8'h8B;
                    16'h109C: data_out = 8'h8C;
                    16'h109D: data_out = 8'h8D;
                    16'h109E: data_out = 8'h8E;
                    16'h109F: data_out = 8'h8F;
                    16'h10A0: data_out = 8'h90;
                    16'h10A1: data_out = 8'h91;
                    16'h10A2: data_out = 8'h92;
                    16'h10A3: data_out = 8'h93;
                    16'h10A4: data_out = 8'h94;
                    16'h10A5: data_out = 8'h95;
                    16'h10A6: data_out = 8'h96;
                    16'h10A7: data_out = 8'h97;
                    16'h10A8: data_out = 8'h98;
                    16'h10A9: data_out = 8'h99;
                    16'h10AA: data_out = 8'h9A;
                    16'h10AB: data_out = 8'h9B;
                    16'h10AC: data_out = 8'h9C;
                    16'h10AD: data_out = 8'h9D;
                    16'h10AE: data_out = 8'h9E;
                    16'h10AF: data_out = 8'h9F;
                    16'h10B0: data_out = 8'hA0;
                    16'h10B1: data_out = 8'hA1;
                    16'h10B2: data_out = 8'hA2;
                    16'h10B3: data_out = 8'hA3;
                    16'h10B4: data_out = 8'hA4;
                    16'h10B5: data_out = 8'hA5;
                    16'h10B6: data_out = 8'hA6;
                    16'h10B7: data_out = 8'hA7;
                    16'h10B8: data_out = 8'hA8;
                    16'h10B9: data_out = 8'hA9;
                    16'h10BA: data_out = 8'hAA;
                    16'h10BB: data_out = 8'hAB;
                    16'h10BC: data_out = 8'hAC;
                    16'h10BD: data_out = 8'hAD;
                    16'h10BE: data_out = 8'hAE;
                    16'h10BF: data_out = 8'hAF;
                    16'h10C0: data_out = 8'hB0;
                    16'h10C1: data_out = 8'hB1;
                    16'h10C2: data_out = 8'hB2;
                    16'h10C3: data_out = 8'hB3;
                    16'h10C4: data_out = 8'hB4;
                    16'h10C5: data_out = 8'hB5;
                    16'h10C6: data_out = 8'hB6;
                    16'h10C7: data_out = 8'hB7;
                    16'h10C8: data_out = 8'hB8;
                    16'h10C9: data_out = 8'hB9;
                    16'h10CA: data_out = 8'hBA;
                    16'h10CB: data_out = 8'hBB;
                    16'h10CC: data_out = 8'hBC;
                    16'h10CD: data_out = 8'hBD;
                    16'h10CE: data_out = 8'hBE;
                    16'h10CF: data_out = 8'hBF;
                    16'h10D0: data_out = 8'hC0;
                    16'h10D1: data_out = 8'hC1;
                    16'h10D2: data_out = 8'hC2;
                    16'h10D3: data_out = 8'hC3;
                    16'h10D4: data_out = 8'hC4;
                    16'h10D5: data_out = 8'hC5;
                    16'h10D6: data_out = 8'hC6;
                    16'h10D7: data_out = 8'hC7;
                    16'h10D8: data_out = 8'hC8;
                    16'h10D9: data_out = 8'hC9;
                    16'h10DA: data_out = 8'hCA;
                    16'h10DB: data_out = 8'hCB;
                    16'h10DC: data_out = 8'hCC;
                    16'h10DD: data_out = 8'hCD;
                    16'h10DE: data_out = 8'hCE;
                    16'h10DF: data_out = 8'hCF;
                    16'h10E0: data_out = 8'hD0;
                    16'h10E1: data_out = 8'hD1;
                    16'h10E2: data_out = 8'hD2;
                    16'h10E3: data_out = 8'hD3;
                    16'h10E4: data_out = 8'hD4;
                    16'h10E5: data_out = 8'hD5;
                    16'h10E6: data_out = 8'hD6;
                    16'h10E7: data_out = 8'hD7;
                    16'h10E8: data_out = 8'hD8;
                    16'h10E9: data_out = 8'hD9;
                    16'h10EA: data_out = 8'hDA;
                    16'h10EB: data_out = 8'hDB;
                    16'h10EC: data_out = 8'hDC;
                    16'h10ED: data_out = 8'hDD;
                    16'h10EE: data_out = 8'hDE;
                    16'h10EF: data_out = 8'hDF;
                    16'h10F0: data_out = 8'hE0;
                    16'h10F1: data_out = 8'hE1;
                    16'h10F2: data_out = 8'hE2;
                    16'h10F3: data_out = 8'hE3;
                    16'h10F4: data_out = 8'hE4;
                    16'h10F5: data_out = 8'hE5;
                    16'h10F6: data_out = 8'hE6;
                    16'h10F7: data_out = 8'hE7;
                    16'h10F8: data_out = 8'hE8;
                    16'h10F9: data_out = 8'hE9;
                    16'h10FA: data_out = 8'hEA;
                    16'h10FB: data_out = 8'hEB;
                    16'h10FC: data_out = 8'hEC;
                    16'h10FD: data_out = 8'hED;
                    16'h10FE: data_out = 8'hEE;
                    16'h10FF: data_out = 8'hEF;
                    16'h1100: data_out = 8'h11;
                    16'h1101: data_out = 8'h12;
                    16'h1102: data_out = 8'h13;
                    16'h1103: data_out = 8'h14;
                    16'h1104: data_out = 8'h15;
                    16'h1105: data_out = 8'h16;
                    16'h1106: data_out = 8'h17;
                    16'h1107: data_out = 8'h18;
                    16'h1108: data_out = 8'h19;
                    16'h1109: data_out = 8'h1A;
                    16'h110A: data_out = 8'h1B;
                    16'h110B: data_out = 8'h1C;
                    16'h110C: data_out = 8'h1D;
                    16'h110D: data_out = 8'h1E;
                    16'h110E: data_out = 8'h1F;
                    16'h110F: data_out = 8'h20;
                    16'h1110: data_out = 8'h21;
                    16'h1111: data_out = 8'h22;
                    16'h1112: data_out = 8'h23;
                    16'h1113: data_out = 8'h24;
                    16'h1114: data_out = 8'h25;
                    16'h1115: data_out = 8'h26;
                    16'h1116: data_out = 8'h27;
                    16'h1117: data_out = 8'h28;
                    16'h1118: data_out = 8'h29;
                    16'h1119: data_out = 8'h2A;
                    16'h111A: data_out = 8'h2B;
                    16'h111B: data_out = 8'h2C;
                    16'h111C: data_out = 8'h2D;
                    16'h111D: data_out = 8'h2E;
                    16'h111E: data_out = 8'h2F;
                    16'h111F: data_out = 8'h30;
                    16'h1120: data_out = 8'h31;
                    16'h1121: data_out = 8'h32;
                    16'h1122: data_out = 8'h33;
                    16'h1123: data_out = 8'h34;
                    16'h1124: data_out = 8'h35;
                    16'h1125: data_out = 8'h36;
                    16'h1126: data_out = 8'h37;
                    16'h1127: data_out = 8'h38;
                    16'h1128: data_out = 8'h39;
                    16'h1129: data_out = 8'h3A;
                    16'h112A: data_out = 8'h3B;
                    16'h112B: data_out = 8'h3C;
                    16'h112C: data_out = 8'h3D;
                    16'h112D: data_out = 8'h3E;
                    16'h112E: data_out = 8'h3F;
                    16'h112F: data_out = 8'h40;
                    16'h1130: data_out = 8'h41;
                    16'h1131: data_out = 8'h42;
                    16'h1132: data_out = 8'h43;
                    16'h1133: data_out = 8'h44;
                    16'h1134: data_out = 8'h45;
                    16'h1135: data_out = 8'h46;
                    16'h1136: data_out = 8'h47;
                    16'h1137: data_out = 8'h48;
                    16'h1138: data_out = 8'h49;
                    16'h1139: data_out = 8'h4A;
                    16'h113A: data_out = 8'h4B;
                    16'h113B: data_out = 8'h4C;
                    16'h113C: data_out = 8'h4D;
                    16'h113D: data_out = 8'h4E;
                    16'h113E: data_out = 8'h4F;
                    16'h113F: data_out = 8'h50;
                    16'h1140: data_out = 8'h51;
                    16'h1141: data_out = 8'h52;
                    16'h1142: data_out = 8'h53;
                    16'h1143: data_out = 8'h54;
                    16'h1144: data_out = 8'h55;
                    16'h1145: data_out = 8'h56;
                    16'h1146: data_out = 8'h57;
                    16'h1147: data_out = 8'h58;
                    16'h1148: data_out = 8'h59;
                    16'h1149: data_out = 8'h5A;
                    16'h114A: data_out = 8'h5B;
                    16'h114B: data_out = 8'h5C;
                    16'h114C: data_out = 8'h5D;
                    16'h114D: data_out = 8'h5E;
                    16'h114E: data_out = 8'h5F;
                    16'h114F: data_out = 8'h60;
                    16'h1150: data_out = 8'h61;
                    16'h1151: data_out = 8'h62;
                    16'h1152: data_out = 8'h63;
                    16'h1153: data_out = 8'h64;
                    16'h1154: data_out = 8'h65;
                    16'h1155: data_out = 8'h66;
                    16'h1156: data_out = 8'h67;
                    16'h1157: data_out = 8'h68;
                    16'h1158: data_out = 8'h69;
                    16'h1159: data_out = 8'h6A;
                    16'h115A: data_out = 8'h6B;
                    16'h115B: data_out = 8'h6C;
                    16'h115C: data_out = 8'h6D;
                    16'h115D: data_out = 8'h6E;
                    16'h115E: data_out = 8'h6F;
                    16'h115F: data_out = 8'h70;
                    16'h1160: data_out = 8'h71;
                    16'h1161: data_out = 8'h72;
                    16'h1162: data_out = 8'h73;
                    16'h1163: data_out = 8'h74;
                    16'h1164: data_out = 8'h75;
                    16'h1165: data_out = 8'h76;
                    16'h1166: data_out = 8'h77;
                    16'h1167: data_out = 8'h78;
                    16'h1168: data_out = 8'h79;
                    16'h1169: data_out = 8'h7A;
                    16'h116A: data_out = 8'h7B;
                    16'h116B: data_out = 8'h7C;
                    16'h116C: data_out = 8'h7D;
                    16'h116D: data_out = 8'h7E;
                    16'h116E: data_out = 8'h7F;
                    16'h116F: data_out = 8'h80;
                    16'h1170: data_out = 8'h81;
                    16'h1171: data_out = 8'h82;
                    16'h1172: data_out = 8'h83;
                    16'h1173: data_out = 8'h84;
                    16'h1174: data_out = 8'h85;
                    16'h1175: data_out = 8'h86;
                    16'h1176: data_out = 8'h87;
                    16'h1177: data_out = 8'h88;
                    16'h1178: data_out = 8'h89;
                    16'h1179: data_out = 8'h8A;
                    16'h117A: data_out = 8'h8B;
                    16'h117B: data_out = 8'h8C;
                    16'h117C: data_out = 8'h8D;
                    16'h117D: data_out = 8'h8E;
                    16'h117E: data_out = 8'h8F;
                    16'h117F: data_out = 8'h90;
                    16'h1180: data_out = 8'h11;
                    16'h1181: data_out = 8'h10;
                    16'h1182: data_out = 8'hF;
                    16'h1183: data_out = 8'hE;
                    16'h1184: data_out = 8'hD;
                    16'h1185: data_out = 8'hC;
                    16'h1186: data_out = 8'hB;
                    16'h1187: data_out = 8'hA;
                    16'h1188: data_out = 8'h9;
                    16'h1189: data_out = 8'h8;
                    16'h118A: data_out = 8'h7;
                    16'h118B: data_out = 8'h6;
                    16'h118C: data_out = 8'h5;
                    16'h118D: data_out = 8'h4;
                    16'h118E: data_out = 8'h3;
                    16'h118F: data_out = 8'h2;
                    16'h1190: data_out = 8'h1;
                    16'h1191: data_out = 8'h0;
                    16'h1192: data_out = 8'h81;
                    16'h1193: data_out = 8'h82;
                    16'h1194: data_out = 8'h83;
                    16'h1195: data_out = 8'h84;
                    16'h1196: data_out = 8'h85;
                    16'h1197: data_out = 8'h86;
                    16'h1198: data_out = 8'h87;
                    16'h1199: data_out = 8'h88;
                    16'h119A: data_out = 8'h89;
                    16'h119B: data_out = 8'h8A;
                    16'h119C: data_out = 8'h8B;
                    16'h119D: data_out = 8'h8C;
                    16'h119E: data_out = 8'h8D;
                    16'h119F: data_out = 8'h8E;
                    16'h11A0: data_out = 8'h8F;
                    16'h11A1: data_out = 8'h90;
                    16'h11A2: data_out = 8'h91;
                    16'h11A3: data_out = 8'h92;
                    16'h11A4: data_out = 8'h93;
                    16'h11A5: data_out = 8'h94;
                    16'h11A6: data_out = 8'h95;
                    16'h11A7: data_out = 8'h96;
                    16'h11A8: data_out = 8'h97;
                    16'h11A9: data_out = 8'h98;
                    16'h11AA: data_out = 8'h99;
                    16'h11AB: data_out = 8'h9A;
                    16'h11AC: data_out = 8'h9B;
                    16'h11AD: data_out = 8'h9C;
                    16'h11AE: data_out = 8'h9D;
                    16'h11AF: data_out = 8'h9E;
                    16'h11B0: data_out = 8'h9F;
                    16'h11B1: data_out = 8'hA0;
                    16'h11B2: data_out = 8'hA1;
                    16'h11B3: data_out = 8'hA2;
                    16'h11B4: data_out = 8'hA3;
                    16'h11B5: data_out = 8'hA4;
                    16'h11B6: data_out = 8'hA5;
                    16'h11B7: data_out = 8'hA6;
                    16'h11B8: data_out = 8'hA7;
                    16'h11B9: data_out = 8'hA8;
                    16'h11BA: data_out = 8'hA9;
                    16'h11BB: data_out = 8'hAA;
                    16'h11BC: data_out = 8'hAB;
                    16'h11BD: data_out = 8'hAC;
                    16'h11BE: data_out = 8'hAD;
                    16'h11BF: data_out = 8'hAE;
                    16'h11C0: data_out = 8'hAF;
                    16'h11C1: data_out = 8'hB0;
                    16'h11C2: data_out = 8'hB1;
                    16'h11C3: data_out = 8'hB2;
                    16'h11C4: data_out = 8'hB3;
                    16'h11C5: data_out = 8'hB4;
                    16'h11C6: data_out = 8'hB5;
                    16'h11C7: data_out = 8'hB6;
                    16'h11C8: data_out = 8'hB7;
                    16'h11C9: data_out = 8'hB8;
                    16'h11CA: data_out = 8'hB9;
                    16'h11CB: data_out = 8'hBA;
                    16'h11CC: data_out = 8'hBB;
                    16'h11CD: data_out = 8'hBC;
                    16'h11CE: data_out = 8'hBD;
                    16'h11CF: data_out = 8'hBE;
                    16'h11D0: data_out = 8'hBF;
                    16'h11D1: data_out = 8'hC0;
                    16'h11D2: data_out = 8'hC1;
                    16'h11D3: data_out = 8'hC2;
                    16'h11D4: data_out = 8'hC3;
                    16'h11D5: data_out = 8'hC4;
                    16'h11D6: data_out = 8'hC5;
                    16'h11D7: data_out = 8'hC6;
                    16'h11D8: data_out = 8'hC7;
                    16'h11D9: data_out = 8'hC8;
                    16'h11DA: data_out = 8'hC9;
                    16'h11DB: data_out = 8'hCA;
                    16'h11DC: data_out = 8'hCB;
                    16'h11DD: data_out = 8'hCC;
                    16'h11DE: data_out = 8'hCD;
                    16'h11DF: data_out = 8'hCE;
                    16'h11E0: data_out = 8'hCF;
                    16'h11E1: data_out = 8'hD0;
                    16'h11E2: data_out = 8'hD1;
                    16'h11E3: data_out = 8'hD2;
                    16'h11E4: data_out = 8'hD3;
                    16'h11E5: data_out = 8'hD4;
                    16'h11E6: data_out = 8'hD5;
                    16'h11E7: data_out = 8'hD6;
                    16'h11E8: data_out = 8'hD7;
                    16'h11E9: data_out = 8'hD8;
                    16'h11EA: data_out = 8'hD9;
                    16'h11EB: data_out = 8'hDA;
                    16'h11EC: data_out = 8'hDB;
                    16'h11ED: data_out = 8'hDC;
                    16'h11EE: data_out = 8'hDD;
                    16'h11EF: data_out = 8'hDE;
                    16'h11F0: data_out = 8'hDF;
                    16'h11F1: data_out = 8'hE0;
                    16'h11F2: data_out = 8'hE1;
                    16'h11F3: data_out = 8'hE2;
                    16'h11F4: data_out = 8'hE3;
                    16'h11F5: data_out = 8'hE4;
                    16'h11F6: data_out = 8'hE5;
                    16'h11F7: data_out = 8'hE6;
                    16'h11F8: data_out = 8'hE7;
                    16'h11F9: data_out = 8'hE8;
                    16'h11FA: data_out = 8'hE9;
                    16'h11FB: data_out = 8'hEA;
                    16'h11FC: data_out = 8'hEB;
                    16'h11FD: data_out = 8'hEC;
                    16'h11FE: data_out = 8'hED;
                    16'h11FF: data_out = 8'hEE;
                    16'h1200: data_out = 8'h12;
                    16'h1201: data_out = 8'h13;
                    16'h1202: data_out = 8'h14;
                    16'h1203: data_out = 8'h15;
                    16'h1204: data_out = 8'h16;
                    16'h1205: data_out = 8'h17;
                    16'h1206: data_out = 8'h18;
                    16'h1207: data_out = 8'h19;
                    16'h1208: data_out = 8'h1A;
                    16'h1209: data_out = 8'h1B;
                    16'h120A: data_out = 8'h1C;
                    16'h120B: data_out = 8'h1D;
                    16'h120C: data_out = 8'h1E;
                    16'h120D: data_out = 8'h1F;
                    16'h120E: data_out = 8'h20;
                    16'h120F: data_out = 8'h21;
                    16'h1210: data_out = 8'h22;
                    16'h1211: data_out = 8'h23;
                    16'h1212: data_out = 8'h24;
                    16'h1213: data_out = 8'h25;
                    16'h1214: data_out = 8'h26;
                    16'h1215: data_out = 8'h27;
                    16'h1216: data_out = 8'h28;
                    16'h1217: data_out = 8'h29;
                    16'h1218: data_out = 8'h2A;
                    16'h1219: data_out = 8'h2B;
                    16'h121A: data_out = 8'h2C;
                    16'h121B: data_out = 8'h2D;
                    16'h121C: data_out = 8'h2E;
                    16'h121D: data_out = 8'h2F;
                    16'h121E: data_out = 8'h30;
                    16'h121F: data_out = 8'h31;
                    16'h1220: data_out = 8'h32;
                    16'h1221: data_out = 8'h33;
                    16'h1222: data_out = 8'h34;
                    16'h1223: data_out = 8'h35;
                    16'h1224: data_out = 8'h36;
                    16'h1225: data_out = 8'h37;
                    16'h1226: data_out = 8'h38;
                    16'h1227: data_out = 8'h39;
                    16'h1228: data_out = 8'h3A;
                    16'h1229: data_out = 8'h3B;
                    16'h122A: data_out = 8'h3C;
                    16'h122B: data_out = 8'h3D;
                    16'h122C: data_out = 8'h3E;
                    16'h122D: data_out = 8'h3F;
                    16'h122E: data_out = 8'h40;
                    16'h122F: data_out = 8'h41;
                    16'h1230: data_out = 8'h42;
                    16'h1231: data_out = 8'h43;
                    16'h1232: data_out = 8'h44;
                    16'h1233: data_out = 8'h45;
                    16'h1234: data_out = 8'h46;
                    16'h1235: data_out = 8'h47;
                    16'h1236: data_out = 8'h48;
                    16'h1237: data_out = 8'h49;
                    16'h1238: data_out = 8'h4A;
                    16'h1239: data_out = 8'h4B;
                    16'h123A: data_out = 8'h4C;
                    16'h123B: data_out = 8'h4D;
                    16'h123C: data_out = 8'h4E;
                    16'h123D: data_out = 8'h4F;
                    16'h123E: data_out = 8'h50;
                    16'h123F: data_out = 8'h51;
                    16'h1240: data_out = 8'h52;
                    16'h1241: data_out = 8'h53;
                    16'h1242: data_out = 8'h54;
                    16'h1243: data_out = 8'h55;
                    16'h1244: data_out = 8'h56;
                    16'h1245: data_out = 8'h57;
                    16'h1246: data_out = 8'h58;
                    16'h1247: data_out = 8'h59;
                    16'h1248: data_out = 8'h5A;
                    16'h1249: data_out = 8'h5B;
                    16'h124A: data_out = 8'h5C;
                    16'h124B: data_out = 8'h5D;
                    16'h124C: data_out = 8'h5E;
                    16'h124D: data_out = 8'h5F;
                    16'h124E: data_out = 8'h60;
                    16'h124F: data_out = 8'h61;
                    16'h1250: data_out = 8'h62;
                    16'h1251: data_out = 8'h63;
                    16'h1252: data_out = 8'h64;
                    16'h1253: data_out = 8'h65;
                    16'h1254: data_out = 8'h66;
                    16'h1255: data_out = 8'h67;
                    16'h1256: data_out = 8'h68;
                    16'h1257: data_out = 8'h69;
                    16'h1258: data_out = 8'h6A;
                    16'h1259: data_out = 8'h6B;
                    16'h125A: data_out = 8'h6C;
                    16'h125B: data_out = 8'h6D;
                    16'h125C: data_out = 8'h6E;
                    16'h125D: data_out = 8'h6F;
                    16'h125E: data_out = 8'h70;
                    16'h125F: data_out = 8'h71;
                    16'h1260: data_out = 8'h72;
                    16'h1261: data_out = 8'h73;
                    16'h1262: data_out = 8'h74;
                    16'h1263: data_out = 8'h75;
                    16'h1264: data_out = 8'h76;
                    16'h1265: data_out = 8'h77;
                    16'h1266: data_out = 8'h78;
                    16'h1267: data_out = 8'h79;
                    16'h1268: data_out = 8'h7A;
                    16'h1269: data_out = 8'h7B;
                    16'h126A: data_out = 8'h7C;
                    16'h126B: data_out = 8'h7D;
                    16'h126C: data_out = 8'h7E;
                    16'h126D: data_out = 8'h7F;
                    16'h126E: data_out = 8'h80;
                    16'h126F: data_out = 8'h81;
                    16'h1270: data_out = 8'h82;
                    16'h1271: data_out = 8'h83;
                    16'h1272: data_out = 8'h84;
                    16'h1273: data_out = 8'h85;
                    16'h1274: data_out = 8'h86;
                    16'h1275: data_out = 8'h87;
                    16'h1276: data_out = 8'h88;
                    16'h1277: data_out = 8'h89;
                    16'h1278: data_out = 8'h8A;
                    16'h1279: data_out = 8'h8B;
                    16'h127A: data_out = 8'h8C;
                    16'h127B: data_out = 8'h8D;
                    16'h127C: data_out = 8'h8E;
                    16'h127D: data_out = 8'h8F;
                    16'h127E: data_out = 8'h90;
                    16'h127F: data_out = 8'h91;
                    16'h1280: data_out = 8'h12;
                    16'h1281: data_out = 8'h11;
                    16'h1282: data_out = 8'h10;
                    16'h1283: data_out = 8'hF;
                    16'h1284: data_out = 8'hE;
                    16'h1285: data_out = 8'hD;
                    16'h1286: data_out = 8'hC;
                    16'h1287: data_out = 8'hB;
                    16'h1288: data_out = 8'hA;
                    16'h1289: data_out = 8'h9;
                    16'h128A: data_out = 8'h8;
                    16'h128B: data_out = 8'h7;
                    16'h128C: data_out = 8'h6;
                    16'h128D: data_out = 8'h5;
                    16'h128E: data_out = 8'h4;
                    16'h128F: data_out = 8'h3;
                    16'h1290: data_out = 8'h2;
                    16'h1291: data_out = 8'h1;
                    16'h1292: data_out = 8'h0;
                    16'h1293: data_out = 8'h81;
                    16'h1294: data_out = 8'h82;
                    16'h1295: data_out = 8'h83;
                    16'h1296: data_out = 8'h84;
                    16'h1297: data_out = 8'h85;
                    16'h1298: data_out = 8'h86;
                    16'h1299: data_out = 8'h87;
                    16'h129A: data_out = 8'h88;
                    16'h129B: data_out = 8'h89;
                    16'h129C: data_out = 8'h8A;
                    16'h129D: data_out = 8'h8B;
                    16'h129E: data_out = 8'h8C;
                    16'h129F: data_out = 8'h8D;
                    16'h12A0: data_out = 8'h8E;
                    16'h12A1: data_out = 8'h8F;
                    16'h12A2: data_out = 8'h90;
                    16'h12A3: data_out = 8'h91;
                    16'h12A4: data_out = 8'h92;
                    16'h12A5: data_out = 8'h93;
                    16'h12A6: data_out = 8'h94;
                    16'h12A7: data_out = 8'h95;
                    16'h12A8: data_out = 8'h96;
                    16'h12A9: data_out = 8'h97;
                    16'h12AA: data_out = 8'h98;
                    16'h12AB: data_out = 8'h99;
                    16'h12AC: data_out = 8'h9A;
                    16'h12AD: data_out = 8'h9B;
                    16'h12AE: data_out = 8'h9C;
                    16'h12AF: data_out = 8'h9D;
                    16'h12B0: data_out = 8'h9E;
                    16'h12B1: data_out = 8'h9F;
                    16'h12B2: data_out = 8'hA0;
                    16'h12B3: data_out = 8'hA1;
                    16'h12B4: data_out = 8'hA2;
                    16'h12B5: data_out = 8'hA3;
                    16'h12B6: data_out = 8'hA4;
                    16'h12B7: data_out = 8'hA5;
                    16'h12B8: data_out = 8'hA6;
                    16'h12B9: data_out = 8'hA7;
                    16'h12BA: data_out = 8'hA8;
                    16'h12BB: data_out = 8'hA9;
                    16'h12BC: data_out = 8'hAA;
                    16'h12BD: data_out = 8'hAB;
                    16'h12BE: data_out = 8'hAC;
                    16'h12BF: data_out = 8'hAD;
                    16'h12C0: data_out = 8'hAE;
                    16'h12C1: data_out = 8'hAF;
                    16'h12C2: data_out = 8'hB0;
                    16'h12C3: data_out = 8'hB1;
                    16'h12C4: data_out = 8'hB2;
                    16'h12C5: data_out = 8'hB3;
                    16'h12C6: data_out = 8'hB4;
                    16'h12C7: data_out = 8'hB5;
                    16'h12C8: data_out = 8'hB6;
                    16'h12C9: data_out = 8'hB7;
                    16'h12CA: data_out = 8'hB8;
                    16'h12CB: data_out = 8'hB9;
                    16'h12CC: data_out = 8'hBA;
                    16'h12CD: data_out = 8'hBB;
                    16'h12CE: data_out = 8'hBC;
                    16'h12CF: data_out = 8'hBD;
                    16'h12D0: data_out = 8'hBE;
                    16'h12D1: data_out = 8'hBF;
                    16'h12D2: data_out = 8'hC0;
                    16'h12D3: data_out = 8'hC1;
                    16'h12D4: data_out = 8'hC2;
                    16'h12D5: data_out = 8'hC3;
                    16'h12D6: data_out = 8'hC4;
                    16'h12D7: data_out = 8'hC5;
                    16'h12D8: data_out = 8'hC6;
                    16'h12D9: data_out = 8'hC7;
                    16'h12DA: data_out = 8'hC8;
                    16'h12DB: data_out = 8'hC9;
                    16'h12DC: data_out = 8'hCA;
                    16'h12DD: data_out = 8'hCB;
                    16'h12DE: data_out = 8'hCC;
                    16'h12DF: data_out = 8'hCD;
                    16'h12E0: data_out = 8'hCE;
                    16'h12E1: data_out = 8'hCF;
                    16'h12E2: data_out = 8'hD0;
                    16'h12E3: data_out = 8'hD1;
                    16'h12E4: data_out = 8'hD2;
                    16'h12E5: data_out = 8'hD3;
                    16'h12E6: data_out = 8'hD4;
                    16'h12E7: data_out = 8'hD5;
                    16'h12E8: data_out = 8'hD6;
                    16'h12E9: data_out = 8'hD7;
                    16'h12EA: data_out = 8'hD8;
                    16'h12EB: data_out = 8'hD9;
                    16'h12EC: data_out = 8'hDA;
                    16'h12ED: data_out = 8'hDB;
                    16'h12EE: data_out = 8'hDC;
                    16'h12EF: data_out = 8'hDD;
                    16'h12F0: data_out = 8'hDE;
                    16'h12F1: data_out = 8'hDF;
                    16'h12F2: data_out = 8'hE0;
                    16'h12F3: data_out = 8'hE1;
                    16'h12F4: data_out = 8'hE2;
                    16'h12F5: data_out = 8'hE3;
                    16'h12F6: data_out = 8'hE4;
                    16'h12F7: data_out = 8'hE5;
                    16'h12F8: data_out = 8'hE6;
                    16'h12F9: data_out = 8'hE7;
                    16'h12FA: data_out = 8'hE8;
                    16'h12FB: data_out = 8'hE9;
                    16'h12FC: data_out = 8'hEA;
                    16'h12FD: data_out = 8'hEB;
                    16'h12FE: data_out = 8'hEC;
                    16'h12FF: data_out = 8'hED;
                    16'h1300: data_out = 8'h13;
                    16'h1301: data_out = 8'h14;
                    16'h1302: data_out = 8'h15;
                    16'h1303: data_out = 8'h16;
                    16'h1304: data_out = 8'h17;
                    16'h1305: data_out = 8'h18;
                    16'h1306: data_out = 8'h19;
                    16'h1307: data_out = 8'h1A;
                    16'h1308: data_out = 8'h1B;
                    16'h1309: data_out = 8'h1C;
                    16'h130A: data_out = 8'h1D;
                    16'h130B: data_out = 8'h1E;
                    16'h130C: data_out = 8'h1F;
                    16'h130D: data_out = 8'h20;
                    16'h130E: data_out = 8'h21;
                    16'h130F: data_out = 8'h22;
                    16'h1310: data_out = 8'h23;
                    16'h1311: data_out = 8'h24;
                    16'h1312: data_out = 8'h25;
                    16'h1313: data_out = 8'h26;
                    16'h1314: data_out = 8'h27;
                    16'h1315: data_out = 8'h28;
                    16'h1316: data_out = 8'h29;
                    16'h1317: data_out = 8'h2A;
                    16'h1318: data_out = 8'h2B;
                    16'h1319: data_out = 8'h2C;
                    16'h131A: data_out = 8'h2D;
                    16'h131B: data_out = 8'h2E;
                    16'h131C: data_out = 8'h2F;
                    16'h131D: data_out = 8'h30;
                    16'h131E: data_out = 8'h31;
                    16'h131F: data_out = 8'h32;
                    16'h1320: data_out = 8'h33;
                    16'h1321: data_out = 8'h34;
                    16'h1322: data_out = 8'h35;
                    16'h1323: data_out = 8'h36;
                    16'h1324: data_out = 8'h37;
                    16'h1325: data_out = 8'h38;
                    16'h1326: data_out = 8'h39;
                    16'h1327: data_out = 8'h3A;
                    16'h1328: data_out = 8'h3B;
                    16'h1329: data_out = 8'h3C;
                    16'h132A: data_out = 8'h3D;
                    16'h132B: data_out = 8'h3E;
                    16'h132C: data_out = 8'h3F;
                    16'h132D: data_out = 8'h40;
                    16'h132E: data_out = 8'h41;
                    16'h132F: data_out = 8'h42;
                    16'h1330: data_out = 8'h43;
                    16'h1331: data_out = 8'h44;
                    16'h1332: data_out = 8'h45;
                    16'h1333: data_out = 8'h46;
                    16'h1334: data_out = 8'h47;
                    16'h1335: data_out = 8'h48;
                    16'h1336: data_out = 8'h49;
                    16'h1337: data_out = 8'h4A;
                    16'h1338: data_out = 8'h4B;
                    16'h1339: data_out = 8'h4C;
                    16'h133A: data_out = 8'h4D;
                    16'h133B: data_out = 8'h4E;
                    16'h133C: data_out = 8'h4F;
                    16'h133D: data_out = 8'h50;
                    16'h133E: data_out = 8'h51;
                    16'h133F: data_out = 8'h52;
                    16'h1340: data_out = 8'h53;
                    16'h1341: data_out = 8'h54;
                    16'h1342: data_out = 8'h55;
                    16'h1343: data_out = 8'h56;
                    16'h1344: data_out = 8'h57;
                    16'h1345: data_out = 8'h58;
                    16'h1346: data_out = 8'h59;
                    16'h1347: data_out = 8'h5A;
                    16'h1348: data_out = 8'h5B;
                    16'h1349: data_out = 8'h5C;
                    16'h134A: data_out = 8'h5D;
                    16'h134B: data_out = 8'h5E;
                    16'h134C: data_out = 8'h5F;
                    16'h134D: data_out = 8'h60;
                    16'h134E: data_out = 8'h61;
                    16'h134F: data_out = 8'h62;
                    16'h1350: data_out = 8'h63;
                    16'h1351: data_out = 8'h64;
                    16'h1352: data_out = 8'h65;
                    16'h1353: data_out = 8'h66;
                    16'h1354: data_out = 8'h67;
                    16'h1355: data_out = 8'h68;
                    16'h1356: data_out = 8'h69;
                    16'h1357: data_out = 8'h6A;
                    16'h1358: data_out = 8'h6B;
                    16'h1359: data_out = 8'h6C;
                    16'h135A: data_out = 8'h6D;
                    16'h135B: data_out = 8'h6E;
                    16'h135C: data_out = 8'h6F;
                    16'h135D: data_out = 8'h70;
                    16'h135E: data_out = 8'h71;
                    16'h135F: data_out = 8'h72;
                    16'h1360: data_out = 8'h73;
                    16'h1361: data_out = 8'h74;
                    16'h1362: data_out = 8'h75;
                    16'h1363: data_out = 8'h76;
                    16'h1364: data_out = 8'h77;
                    16'h1365: data_out = 8'h78;
                    16'h1366: data_out = 8'h79;
                    16'h1367: data_out = 8'h7A;
                    16'h1368: data_out = 8'h7B;
                    16'h1369: data_out = 8'h7C;
                    16'h136A: data_out = 8'h7D;
                    16'h136B: data_out = 8'h7E;
                    16'h136C: data_out = 8'h7F;
                    16'h136D: data_out = 8'h80;
                    16'h136E: data_out = 8'h81;
                    16'h136F: data_out = 8'h82;
                    16'h1370: data_out = 8'h83;
                    16'h1371: data_out = 8'h84;
                    16'h1372: data_out = 8'h85;
                    16'h1373: data_out = 8'h86;
                    16'h1374: data_out = 8'h87;
                    16'h1375: data_out = 8'h88;
                    16'h1376: data_out = 8'h89;
                    16'h1377: data_out = 8'h8A;
                    16'h1378: data_out = 8'h8B;
                    16'h1379: data_out = 8'h8C;
                    16'h137A: data_out = 8'h8D;
                    16'h137B: data_out = 8'h8E;
                    16'h137C: data_out = 8'h8F;
                    16'h137D: data_out = 8'h90;
                    16'h137E: data_out = 8'h91;
                    16'h137F: data_out = 8'h92;
                    16'h1380: data_out = 8'h13;
                    16'h1381: data_out = 8'h12;
                    16'h1382: data_out = 8'h11;
                    16'h1383: data_out = 8'h10;
                    16'h1384: data_out = 8'hF;
                    16'h1385: data_out = 8'hE;
                    16'h1386: data_out = 8'hD;
                    16'h1387: data_out = 8'hC;
                    16'h1388: data_out = 8'hB;
                    16'h1389: data_out = 8'hA;
                    16'h138A: data_out = 8'h9;
                    16'h138B: data_out = 8'h8;
                    16'h138C: data_out = 8'h7;
                    16'h138D: data_out = 8'h6;
                    16'h138E: data_out = 8'h5;
                    16'h138F: data_out = 8'h4;
                    16'h1390: data_out = 8'h3;
                    16'h1391: data_out = 8'h2;
                    16'h1392: data_out = 8'h1;
                    16'h1393: data_out = 8'h0;
                    16'h1394: data_out = 8'h81;
                    16'h1395: data_out = 8'h82;
                    16'h1396: data_out = 8'h83;
                    16'h1397: data_out = 8'h84;
                    16'h1398: data_out = 8'h85;
                    16'h1399: data_out = 8'h86;
                    16'h139A: data_out = 8'h87;
                    16'h139B: data_out = 8'h88;
                    16'h139C: data_out = 8'h89;
                    16'h139D: data_out = 8'h8A;
                    16'h139E: data_out = 8'h8B;
                    16'h139F: data_out = 8'h8C;
                    16'h13A0: data_out = 8'h8D;
                    16'h13A1: data_out = 8'h8E;
                    16'h13A2: data_out = 8'h8F;
                    16'h13A3: data_out = 8'h90;
                    16'h13A4: data_out = 8'h91;
                    16'h13A5: data_out = 8'h92;
                    16'h13A6: data_out = 8'h93;
                    16'h13A7: data_out = 8'h94;
                    16'h13A8: data_out = 8'h95;
                    16'h13A9: data_out = 8'h96;
                    16'h13AA: data_out = 8'h97;
                    16'h13AB: data_out = 8'h98;
                    16'h13AC: data_out = 8'h99;
                    16'h13AD: data_out = 8'h9A;
                    16'h13AE: data_out = 8'h9B;
                    16'h13AF: data_out = 8'h9C;
                    16'h13B0: data_out = 8'h9D;
                    16'h13B1: data_out = 8'h9E;
                    16'h13B2: data_out = 8'h9F;
                    16'h13B3: data_out = 8'hA0;
                    16'h13B4: data_out = 8'hA1;
                    16'h13B5: data_out = 8'hA2;
                    16'h13B6: data_out = 8'hA3;
                    16'h13B7: data_out = 8'hA4;
                    16'h13B8: data_out = 8'hA5;
                    16'h13B9: data_out = 8'hA6;
                    16'h13BA: data_out = 8'hA7;
                    16'h13BB: data_out = 8'hA8;
                    16'h13BC: data_out = 8'hA9;
                    16'h13BD: data_out = 8'hAA;
                    16'h13BE: data_out = 8'hAB;
                    16'h13BF: data_out = 8'hAC;
                    16'h13C0: data_out = 8'hAD;
                    16'h13C1: data_out = 8'hAE;
                    16'h13C2: data_out = 8'hAF;
                    16'h13C3: data_out = 8'hB0;
                    16'h13C4: data_out = 8'hB1;
                    16'h13C5: data_out = 8'hB2;
                    16'h13C6: data_out = 8'hB3;
                    16'h13C7: data_out = 8'hB4;
                    16'h13C8: data_out = 8'hB5;
                    16'h13C9: data_out = 8'hB6;
                    16'h13CA: data_out = 8'hB7;
                    16'h13CB: data_out = 8'hB8;
                    16'h13CC: data_out = 8'hB9;
                    16'h13CD: data_out = 8'hBA;
                    16'h13CE: data_out = 8'hBB;
                    16'h13CF: data_out = 8'hBC;
                    16'h13D0: data_out = 8'hBD;
                    16'h13D1: data_out = 8'hBE;
                    16'h13D2: data_out = 8'hBF;
                    16'h13D3: data_out = 8'hC0;
                    16'h13D4: data_out = 8'hC1;
                    16'h13D5: data_out = 8'hC2;
                    16'h13D6: data_out = 8'hC3;
                    16'h13D7: data_out = 8'hC4;
                    16'h13D8: data_out = 8'hC5;
                    16'h13D9: data_out = 8'hC6;
                    16'h13DA: data_out = 8'hC7;
                    16'h13DB: data_out = 8'hC8;
                    16'h13DC: data_out = 8'hC9;
                    16'h13DD: data_out = 8'hCA;
                    16'h13DE: data_out = 8'hCB;
                    16'h13DF: data_out = 8'hCC;
                    16'h13E0: data_out = 8'hCD;
                    16'h13E1: data_out = 8'hCE;
                    16'h13E2: data_out = 8'hCF;
                    16'h13E3: data_out = 8'hD0;
                    16'h13E4: data_out = 8'hD1;
                    16'h13E5: data_out = 8'hD2;
                    16'h13E6: data_out = 8'hD3;
                    16'h13E7: data_out = 8'hD4;
                    16'h13E8: data_out = 8'hD5;
                    16'h13E9: data_out = 8'hD6;
                    16'h13EA: data_out = 8'hD7;
                    16'h13EB: data_out = 8'hD8;
                    16'h13EC: data_out = 8'hD9;
                    16'h13ED: data_out = 8'hDA;
                    16'h13EE: data_out = 8'hDB;
                    16'h13EF: data_out = 8'hDC;
                    16'h13F0: data_out = 8'hDD;
                    16'h13F1: data_out = 8'hDE;
                    16'h13F2: data_out = 8'hDF;
                    16'h13F3: data_out = 8'hE0;
                    16'h13F4: data_out = 8'hE1;
                    16'h13F5: data_out = 8'hE2;
                    16'h13F6: data_out = 8'hE3;
                    16'h13F7: data_out = 8'hE4;
                    16'h13F8: data_out = 8'hE5;
                    16'h13F9: data_out = 8'hE6;
                    16'h13FA: data_out = 8'hE7;
                    16'h13FB: data_out = 8'hE8;
                    16'h13FC: data_out = 8'hE9;
                    16'h13FD: data_out = 8'hEA;
                    16'h13FE: data_out = 8'hEB;
                    16'h13FF: data_out = 8'hEC;
                    16'h1400: data_out = 8'h14;
                    16'h1401: data_out = 8'h15;
                    16'h1402: data_out = 8'h16;
                    16'h1403: data_out = 8'h17;
                    16'h1404: data_out = 8'h18;
                    16'h1405: data_out = 8'h19;
                    16'h1406: data_out = 8'h1A;
                    16'h1407: data_out = 8'h1B;
                    16'h1408: data_out = 8'h1C;
                    16'h1409: data_out = 8'h1D;
                    16'h140A: data_out = 8'h1E;
                    16'h140B: data_out = 8'h1F;
                    16'h140C: data_out = 8'h20;
                    16'h140D: data_out = 8'h21;
                    16'h140E: data_out = 8'h22;
                    16'h140F: data_out = 8'h23;
                    16'h1410: data_out = 8'h24;
                    16'h1411: data_out = 8'h25;
                    16'h1412: data_out = 8'h26;
                    16'h1413: data_out = 8'h27;
                    16'h1414: data_out = 8'h28;
                    16'h1415: data_out = 8'h29;
                    16'h1416: data_out = 8'h2A;
                    16'h1417: data_out = 8'h2B;
                    16'h1418: data_out = 8'h2C;
                    16'h1419: data_out = 8'h2D;
                    16'h141A: data_out = 8'h2E;
                    16'h141B: data_out = 8'h2F;
                    16'h141C: data_out = 8'h30;
                    16'h141D: data_out = 8'h31;
                    16'h141E: data_out = 8'h32;
                    16'h141F: data_out = 8'h33;
                    16'h1420: data_out = 8'h34;
                    16'h1421: data_out = 8'h35;
                    16'h1422: data_out = 8'h36;
                    16'h1423: data_out = 8'h37;
                    16'h1424: data_out = 8'h38;
                    16'h1425: data_out = 8'h39;
                    16'h1426: data_out = 8'h3A;
                    16'h1427: data_out = 8'h3B;
                    16'h1428: data_out = 8'h3C;
                    16'h1429: data_out = 8'h3D;
                    16'h142A: data_out = 8'h3E;
                    16'h142B: data_out = 8'h3F;
                    16'h142C: data_out = 8'h40;
                    16'h142D: data_out = 8'h41;
                    16'h142E: data_out = 8'h42;
                    16'h142F: data_out = 8'h43;
                    16'h1430: data_out = 8'h44;
                    16'h1431: data_out = 8'h45;
                    16'h1432: data_out = 8'h46;
                    16'h1433: data_out = 8'h47;
                    16'h1434: data_out = 8'h48;
                    16'h1435: data_out = 8'h49;
                    16'h1436: data_out = 8'h4A;
                    16'h1437: data_out = 8'h4B;
                    16'h1438: data_out = 8'h4C;
                    16'h1439: data_out = 8'h4D;
                    16'h143A: data_out = 8'h4E;
                    16'h143B: data_out = 8'h4F;
                    16'h143C: data_out = 8'h50;
                    16'h143D: data_out = 8'h51;
                    16'h143E: data_out = 8'h52;
                    16'h143F: data_out = 8'h53;
                    16'h1440: data_out = 8'h54;
                    16'h1441: data_out = 8'h55;
                    16'h1442: data_out = 8'h56;
                    16'h1443: data_out = 8'h57;
                    16'h1444: data_out = 8'h58;
                    16'h1445: data_out = 8'h59;
                    16'h1446: data_out = 8'h5A;
                    16'h1447: data_out = 8'h5B;
                    16'h1448: data_out = 8'h5C;
                    16'h1449: data_out = 8'h5D;
                    16'h144A: data_out = 8'h5E;
                    16'h144B: data_out = 8'h5F;
                    16'h144C: data_out = 8'h60;
                    16'h144D: data_out = 8'h61;
                    16'h144E: data_out = 8'h62;
                    16'h144F: data_out = 8'h63;
                    16'h1450: data_out = 8'h64;
                    16'h1451: data_out = 8'h65;
                    16'h1452: data_out = 8'h66;
                    16'h1453: data_out = 8'h67;
                    16'h1454: data_out = 8'h68;
                    16'h1455: data_out = 8'h69;
                    16'h1456: data_out = 8'h6A;
                    16'h1457: data_out = 8'h6B;
                    16'h1458: data_out = 8'h6C;
                    16'h1459: data_out = 8'h6D;
                    16'h145A: data_out = 8'h6E;
                    16'h145B: data_out = 8'h6F;
                    16'h145C: data_out = 8'h70;
                    16'h145D: data_out = 8'h71;
                    16'h145E: data_out = 8'h72;
                    16'h145F: data_out = 8'h73;
                    16'h1460: data_out = 8'h74;
                    16'h1461: data_out = 8'h75;
                    16'h1462: data_out = 8'h76;
                    16'h1463: data_out = 8'h77;
                    16'h1464: data_out = 8'h78;
                    16'h1465: data_out = 8'h79;
                    16'h1466: data_out = 8'h7A;
                    16'h1467: data_out = 8'h7B;
                    16'h1468: data_out = 8'h7C;
                    16'h1469: data_out = 8'h7D;
                    16'h146A: data_out = 8'h7E;
                    16'h146B: data_out = 8'h7F;
                    16'h146C: data_out = 8'h80;
                    16'h146D: data_out = 8'h81;
                    16'h146E: data_out = 8'h82;
                    16'h146F: data_out = 8'h83;
                    16'h1470: data_out = 8'h84;
                    16'h1471: data_out = 8'h85;
                    16'h1472: data_out = 8'h86;
                    16'h1473: data_out = 8'h87;
                    16'h1474: data_out = 8'h88;
                    16'h1475: data_out = 8'h89;
                    16'h1476: data_out = 8'h8A;
                    16'h1477: data_out = 8'h8B;
                    16'h1478: data_out = 8'h8C;
                    16'h1479: data_out = 8'h8D;
                    16'h147A: data_out = 8'h8E;
                    16'h147B: data_out = 8'h8F;
                    16'h147C: data_out = 8'h90;
                    16'h147D: data_out = 8'h91;
                    16'h147E: data_out = 8'h92;
                    16'h147F: data_out = 8'h93;
                    16'h1480: data_out = 8'h14;
                    16'h1481: data_out = 8'h13;
                    16'h1482: data_out = 8'h12;
                    16'h1483: data_out = 8'h11;
                    16'h1484: data_out = 8'h10;
                    16'h1485: data_out = 8'hF;
                    16'h1486: data_out = 8'hE;
                    16'h1487: data_out = 8'hD;
                    16'h1488: data_out = 8'hC;
                    16'h1489: data_out = 8'hB;
                    16'h148A: data_out = 8'hA;
                    16'h148B: data_out = 8'h9;
                    16'h148C: data_out = 8'h8;
                    16'h148D: data_out = 8'h7;
                    16'h148E: data_out = 8'h6;
                    16'h148F: data_out = 8'h5;
                    16'h1490: data_out = 8'h4;
                    16'h1491: data_out = 8'h3;
                    16'h1492: data_out = 8'h2;
                    16'h1493: data_out = 8'h1;
                    16'h1494: data_out = 8'h0;
                    16'h1495: data_out = 8'h81;
                    16'h1496: data_out = 8'h82;
                    16'h1497: data_out = 8'h83;
                    16'h1498: data_out = 8'h84;
                    16'h1499: data_out = 8'h85;
                    16'h149A: data_out = 8'h86;
                    16'h149B: data_out = 8'h87;
                    16'h149C: data_out = 8'h88;
                    16'h149D: data_out = 8'h89;
                    16'h149E: data_out = 8'h8A;
                    16'h149F: data_out = 8'h8B;
                    16'h14A0: data_out = 8'h8C;
                    16'h14A1: data_out = 8'h8D;
                    16'h14A2: data_out = 8'h8E;
                    16'h14A3: data_out = 8'h8F;
                    16'h14A4: data_out = 8'h90;
                    16'h14A5: data_out = 8'h91;
                    16'h14A6: data_out = 8'h92;
                    16'h14A7: data_out = 8'h93;
                    16'h14A8: data_out = 8'h94;
                    16'h14A9: data_out = 8'h95;
                    16'h14AA: data_out = 8'h96;
                    16'h14AB: data_out = 8'h97;
                    16'h14AC: data_out = 8'h98;
                    16'h14AD: data_out = 8'h99;
                    16'h14AE: data_out = 8'h9A;
                    16'h14AF: data_out = 8'h9B;
                    16'h14B0: data_out = 8'h9C;
                    16'h14B1: data_out = 8'h9D;
                    16'h14B2: data_out = 8'h9E;
                    16'h14B3: data_out = 8'h9F;
                    16'h14B4: data_out = 8'hA0;
                    16'h14B5: data_out = 8'hA1;
                    16'h14B6: data_out = 8'hA2;
                    16'h14B7: data_out = 8'hA3;
                    16'h14B8: data_out = 8'hA4;
                    16'h14B9: data_out = 8'hA5;
                    16'h14BA: data_out = 8'hA6;
                    16'h14BB: data_out = 8'hA7;
                    16'h14BC: data_out = 8'hA8;
                    16'h14BD: data_out = 8'hA9;
                    16'h14BE: data_out = 8'hAA;
                    16'h14BF: data_out = 8'hAB;
                    16'h14C0: data_out = 8'hAC;
                    16'h14C1: data_out = 8'hAD;
                    16'h14C2: data_out = 8'hAE;
                    16'h14C3: data_out = 8'hAF;
                    16'h14C4: data_out = 8'hB0;
                    16'h14C5: data_out = 8'hB1;
                    16'h14C6: data_out = 8'hB2;
                    16'h14C7: data_out = 8'hB3;
                    16'h14C8: data_out = 8'hB4;
                    16'h14C9: data_out = 8'hB5;
                    16'h14CA: data_out = 8'hB6;
                    16'h14CB: data_out = 8'hB7;
                    16'h14CC: data_out = 8'hB8;
                    16'h14CD: data_out = 8'hB9;
                    16'h14CE: data_out = 8'hBA;
                    16'h14CF: data_out = 8'hBB;
                    16'h14D0: data_out = 8'hBC;
                    16'h14D1: data_out = 8'hBD;
                    16'h14D2: data_out = 8'hBE;
                    16'h14D3: data_out = 8'hBF;
                    16'h14D4: data_out = 8'hC0;
                    16'h14D5: data_out = 8'hC1;
                    16'h14D6: data_out = 8'hC2;
                    16'h14D7: data_out = 8'hC3;
                    16'h14D8: data_out = 8'hC4;
                    16'h14D9: data_out = 8'hC5;
                    16'h14DA: data_out = 8'hC6;
                    16'h14DB: data_out = 8'hC7;
                    16'h14DC: data_out = 8'hC8;
                    16'h14DD: data_out = 8'hC9;
                    16'h14DE: data_out = 8'hCA;
                    16'h14DF: data_out = 8'hCB;
                    16'h14E0: data_out = 8'hCC;
                    16'h14E1: data_out = 8'hCD;
                    16'h14E2: data_out = 8'hCE;
                    16'h14E3: data_out = 8'hCF;
                    16'h14E4: data_out = 8'hD0;
                    16'h14E5: data_out = 8'hD1;
                    16'h14E6: data_out = 8'hD2;
                    16'h14E7: data_out = 8'hD3;
                    16'h14E8: data_out = 8'hD4;
                    16'h14E9: data_out = 8'hD5;
                    16'h14EA: data_out = 8'hD6;
                    16'h14EB: data_out = 8'hD7;
                    16'h14EC: data_out = 8'hD8;
                    16'h14ED: data_out = 8'hD9;
                    16'h14EE: data_out = 8'hDA;
                    16'h14EF: data_out = 8'hDB;
                    16'h14F0: data_out = 8'hDC;
                    16'h14F1: data_out = 8'hDD;
                    16'h14F2: data_out = 8'hDE;
                    16'h14F3: data_out = 8'hDF;
                    16'h14F4: data_out = 8'hE0;
                    16'h14F5: data_out = 8'hE1;
                    16'h14F6: data_out = 8'hE2;
                    16'h14F7: data_out = 8'hE3;
                    16'h14F8: data_out = 8'hE4;
                    16'h14F9: data_out = 8'hE5;
                    16'h14FA: data_out = 8'hE6;
                    16'h14FB: data_out = 8'hE7;
                    16'h14FC: data_out = 8'hE8;
                    16'h14FD: data_out = 8'hE9;
                    16'h14FE: data_out = 8'hEA;
                    16'h14FF: data_out = 8'hEB;
                    16'h1500: data_out = 8'h15;
                    16'h1501: data_out = 8'h16;
                    16'h1502: data_out = 8'h17;
                    16'h1503: data_out = 8'h18;
                    16'h1504: data_out = 8'h19;
                    16'h1505: data_out = 8'h1A;
                    16'h1506: data_out = 8'h1B;
                    16'h1507: data_out = 8'h1C;
                    16'h1508: data_out = 8'h1D;
                    16'h1509: data_out = 8'h1E;
                    16'h150A: data_out = 8'h1F;
                    16'h150B: data_out = 8'h20;
                    16'h150C: data_out = 8'h21;
                    16'h150D: data_out = 8'h22;
                    16'h150E: data_out = 8'h23;
                    16'h150F: data_out = 8'h24;
                    16'h1510: data_out = 8'h25;
                    16'h1511: data_out = 8'h26;
                    16'h1512: data_out = 8'h27;
                    16'h1513: data_out = 8'h28;
                    16'h1514: data_out = 8'h29;
                    16'h1515: data_out = 8'h2A;
                    16'h1516: data_out = 8'h2B;
                    16'h1517: data_out = 8'h2C;
                    16'h1518: data_out = 8'h2D;
                    16'h1519: data_out = 8'h2E;
                    16'h151A: data_out = 8'h2F;
                    16'h151B: data_out = 8'h30;
                    16'h151C: data_out = 8'h31;
                    16'h151D: data_out = 8'h32;
                    16'h151E: data_out = 8'h33;
                    16'h151F: data_out = 8'h34;
                    16'h1520: data_out = 8'h35;
                    16'h1521: data_out = 8'h36;
                    16'h1522: data_out = 8'h37;
                    16'h1523: data_out = 8'h38;
                    16'h1524: data_out = 8'h39;
                    16'h1525: data_out = 8'h3A;
                    16'h1526: data_out = 8'h3B;
                    16'h1527: data_out = 8'h3C;
                    16'h1528: data_out = 8'h3D;
                    16'h1529: data_out = 8'h3E;
                    16'h152A: data_out = 8'h3F;
                    16'h152B: data_out = 8'h40;
                    16'h152C: data_out = 8'h41;
                    16'h152D: data_out = 8'h42;
                    16'h152E: data_out = 8'h43;
                    16'h152F: data_out = 8'h44;
                    16'h1530: data_out = 8'h45;
                    16'h1531: data_out = 8'h46;
                    16'h1532: data_out = 8'h47;
                    16'h1533: data_out = 8'h48;
                    16'h1534: data_out = 8'h49;
                    16'h1535: data_out = 8'h4A;
                    16'h1536: data_out = 8'h4B;
                    16'h1537: data_out = 8'h4C;
                    16'h1538: data_out = 8'h4D;
                    16'h1539: data_out = 8'h4E;
                    16'h153A: data_out = 8'h4F;
                    16'h153B: data_out = 8'h50;
                    16'h153C: data_out = 8'h51;
                    16'h153D: data_out = 8'h52;
                    16'h153E: data_out = 8'h53;
                    16'h153F: data_out = 8'h54;
                    16'h1540: data_out = 8'h55;
                    16'h1541: data_out = 8'h56;
                    16'h1542: data_out = 8'h57;
                    16'h1543: data_out = 8'h58;
                    16'h1544: data_out = 8'h59;
                    16'h1545: data_out = 8'h5A;
                    16'h1546: data_out = 8'h5B;
                    16'h1547: data_out = 8'h5C;
                    16'h1548: data_out = 8'h5D;
                    16'h1549: data_out = 8'h5E;
                    16'h154A: data_out = 8'h5F;
                    16'h154B: data_out = 8'h60;
                    16'h154C: data_out = 8'h61;
                    16'h154D: data_out = 8'h62;
                    16'h154E: data_out = 8'h63;
                    16'h154F: data_out = 8'h64;
                    16'h1550: data_out = 8'h65;
                    16'h1551: data_out = 8'h66;
                    16'h1552: data_out = 8'h67;
                    16'h1553: data_out = 8'h68;
                    16'h1554: data_out = 8'h69;
                    16'h1555: data_out = 8'h6A;
                    16'h1556: data_out = 8'h6B;
                    16'h1557: data_out = 8'h6C;
                    16'h1558: data_out = 8'h6D;
                    16'h1559: data_out = 8'h6E;
                    16'h155A: data_out = 8'h6F;
                    16'h155B: data_out = 8'h70;
                    16'h155C: data_out = 8'h71;
                    16'h155D: data_out = 8'h72;
                    16'h155E: data_out = 8'h73;
                    16'h155F: data_out = 8'h74;
                    16'h1560: data_out = 8'h75;
                    16'h1561: data_out = 8'h76;
                    16'h1562: data_out = 8'h77;
                    16'h1563: data_out = 8'h78;
                    16'h1564: data_out = 8'h79;
                    16'h1565: data_out = 8'h7A;
                    16'h1566: data_out = 8'h7B;
                    16'h1567: data_out = 8'h7C;
                    16'h1568: data_out = 8'h7D;
                    16'h1569: data_out = 8'h7E;
                    16'h156A: data_out = 8'h7F;
                    16'h156B: data_out = 8'h80;
                    16'h156C: data_out = 8'h81;
                    16'h156D: data_out = 8'h82;
                    16'h156E: data_out = 8'h83;
                    16'h156F: data_out = 8'h84;
                    16'h1570: data_out = 8'h85;
                    16'h1571: data_out = 8'h86;
                    16'h1572: data_out = 8'h87;
                    16'h1573: data_out = 8'h88;
                    16'h1574: data_out = 8'h89;
                    16'h1575: data_out = 8'h8A;
                    16'h1576: data_out = 8'h8B;
                    16'h1577: data_out = 8'h8C;
                    16'h1578: data_out = 8'h8D;
                    16'h1579: data_out = 8'h8E;
                    16'h157A: data_out = 8'h8F;
                    16'h157B: data_out = 8'h90;
                    16'h157C: data_out = 8'h91;
                    16'h157D: data_out = 8'h92;
                    16'h157E: data_out = 8'h93;
                    16'h157F: data_out = 8'h94;
                    16'h1580: data_out = 8'h15;
                    16'h1581: data_out = 8'h14;
                    16'h1582: data_out = 8'h13;
                    16'h1583: data_out = 8'h12;
                    16'h1584: data_out = 8'h11;
                    16'h1585: data_out = 8'h10;
                    16'h1586: data_out = 8'hF;
                    16'h1587: data_out = 8'hE;
                    16'h1588: data_out = 8'hD;
                    16'h1589: data_out = 8'hC;
                    16'h158A: data_out = 8'hB;
                    16'h158B: data_out = 8'hA;
                    16'h158C: data_out = 8'h9;
                    16'h158D: data_out = 8'h8;
                    16'h158E: data_out = 8'h7;
                    16'h158F: data_out = 8'h6;
                    16'h1590: data_out = 8'h5;
                    16'h1591: data_out = 8'h4;
                    16'h1592: data_out = 8'h3;
                    16'h1593: data_out = 8'h2;
                    16'h1594: data_out = 8'h1;
                    16'h1595: data_out = 8'h0;
                    16'h1596: data_out = 8'h81;
                    16'h1597: data_out = 8'h82;
                    16'h1598: data_out = 8'h83;
                    16'h1599: data_out = 8'h84;
                    16'h159A: data_out = 8'h85;
                    16'h159B: data_out = 8'h86;
                    16'h159C: data_out = 8'h87;
                    16'h159D: data_out = 8'h88;
                    16'h159E: data_out = 8'h89;
                    16'h159F: data_out = 8'h8A;
                    16'h15A0: data_out = 8'h8B;
                    16'h15A1: data_out = 8'h8C;
                    16'h15A2: data_out = 8'h8D;
                    16'h15A3: data_out = 8'h8E;
                    16'h15A4: data_out = 8'h8F;
                    16'h15A5: data_out = 8'h90;
                    16'h15A6: data_out = 8'h91;
                    16'h15A7: data_out = 8'h92;
                    16'h15A8: data_out = 8'h93;
                    16'h15A9: data_out = 8'h94;
                    16'h15AA: data_out = 8'h95;
                    16'h15AB: data_out = 8'h96;
                    16'h15AC: data_out = 8'h97;
                    16'h15AD: data_out = 8'h98;
                    16'h15AE: data_out = 8'h99;
                    16'h15AF: data_out = 8'h9A;
                    16'h15B0: data_out = 8'h9B;
                    16'h15B1: data_out = 8'h9C;
                    16'h15B2: data_out = 8'h9D;
                    16'h15B3: data_out = 8'h9E;
                    16'h15B4: data_out = 8'h9F;
                    16'h15B5: data_out = 8'hA0;
                    16'h15B6: data_out = 8'hA1;
                    16'h15B7: data_out = 8'hA2;
                    16'h15B8: data_out = 8'hA3;
                    16'h15B9: data_out = 8'hA4;
                    16'h15BA: data_out = 8'hA5;
                    16'h15BB: data_out = 8'hA6;
                    16'h15BC: data_out = 8'hA7;
                    16'h15BD: data_out = 8'hA8;
                    16'h15BE: data_out = 8'hA9;
                    16'h15BF: data_out = 8'hAA;
                    16'h15C0: data_out = 8'hAB;
                    16'h15C1: data_out = 8'hAC;
                    16'h15C2: data_out = 8'hAD;
                    16'h15C3: data_out = 8'hAE;
                    16'h15C4: data_out = 8'hAF;
                    16'h15C5: data_out = 8'hB0;
                    16'h15C6: data_out = 8'hB1;
                    16'h15C7: data_out = 8'hB2;
                    16'h15C8: data_out = 8'hB3;
                    16'h15C9: data_out = 8'hB4;
                    16'h15CA: data_out = 8'hB5;
                    16'h15CB: data_out = 8'hB6;
                    16'h15CC: data_out = 8'hB7;
                    16'h15CD: data_out = 8'hB8;
                    16'h15CE: data_out = 8'hB9;
                    16'h15CF: data_out = 8'hBA;
                    16'h15D0: data_out = 8'hBB;
                    16'h15D1: data_out = 8'hBC;
                    16'h15D2: data_out = 8'hBD;
                    16'h15D3: data_out = 8'hBE;
                    16'h15D4: data_out = 8'hBF;
                    16'h15D5: data_out = 8'hC0;
                    16'h15D6: data_out = 8'hC1;
                    16'h15D7: data_out = 8'hC2;
                    16'h15D8: data_out = 8'hC3;
                    16'h15D9: data_out = 8'hC4;
                    16'h15DA: data_out = 8'hC5;
                    16'h15DB: data_out = 8'hC6;
                    16'h15DC: data_out = 8'hC7;
                    16'h15DD: data_out = 8'hC8;
                    16'h15DE: data_out = 8'hC9;
                    16'h15DF: data_out = 8'hCA;
                    16'h15E0: data_out = 8'hCB;
                    16'h15E1: data_out = 8'hCC;
                    16'h15E2: data_out = 8'hCD;
                    16'h15E3: data_out = 8'hCE;
                    16'h15E4: data_out = 8'hCF;
                    16'h15E5: data_out = 8'hD0;
                    16'h15E6: data_out = 8'hD1;
                    16'h15E7: data_out = 8'hD2;
                    16'h15E8: data_out = 8'hD3;
                    16'h15E9: data_out = 8'hD4;
                    16'h15EA: data_out = 8'hD5;
                    16'h15EB: data_out = 8'hD6;
                    16'h15EC: data_out = 8'hD7;
                    16'h15ED: data_out = 8'hD8;
                    16'h15EE: data_out = 8'hD9;
                    16'h15EF: data_out = 8'hDA;
                    16'h15F0: data_out = 8'hDB;
                    16'h15F1: data_out = 8'hDC;
                    16'h15F2: data_out = 8'hDD;
                    16'h15F3: data_out = 8'hDE;
                    16'h15F4: data_out = 8'hDF;
                    16'h15F5: data_out = 8'hE0;
                    16'h15F6: data_out = 8'hE1;
                    16'h15F7: data_out = 8'hE2;
                    16'h15F8: data_out = 8'hE3;
                    16'h15F9: data_out = 8'hE4;
                    16'h15FA: data_out = 8'hE5;
                    16'h15FB: data_out = 8'hE6;
                    16'h15FC: data_out = 8'hE7;
                    16'h15FD: data_out = 8'hE8;
                    16'h15FE: data_out = 8'hE9;
                    16'h15FF: data_out = 8'hEA;
                    16'h1600: data_out = 8'h16;
                    16'h1601: data_out = 8'h17;
                    16'h1602: data_out = 8'h18;
                    16'h1603: data_out = 8'h19;
                    16'h1604: data_out = 8'h1A;
                    16'h1605: data_out = 8'h1B;
                    16'h1606: data_out = 8'h1C;
                    16'h1607: data_out = 8'h1D;
                    16'h1608: data_out = 8'h1E;
                    16'h1609: data_out = 8'h1F;
                    16'h160A: data_out = 8'h20;
                    16'h160B: data_out = 8'h21;
                    16'h160C: data_out = 8'h22;
                    16'h160D: data_out = 8'h23;
                    16'h160E: data_out = 8'h24;
                    16'h160F: data_out = 8'h25;
                    16'h1610: data_out = 8'h26;
                    16'h1611: data_out = 8'h27;
                    16'h1612: data_out = 8'h28;
                    16'h1613: data_out = 8'h29;
                    16'h1614: data_out = 8'h2A;
                    16'h1615: data_out = 8'h2B;
                    16'h1616: data_out = 8'h2C;
                    16'h1617: data_out = 8'h2D;
                    16'h1618: data_out = 8'h2E;
                    16'h1619: data_out = 8'h2F;
                    16'h161A: data_out = 8'h30;
                    16'h161B: data_out = 8'h31;
                    16'h161C: data_out = 8'h32;
                    16'h161D: data_out = 8'h33;
                    16'h161E: data_out = 8'h34;
                    16'h161F: data_out = 8'h35;
                    16'h1620: data_out = 8'h36;
                    16'h1621: data_out = 8'h37;
                    16'h1622: data_out = 8'h38;
                    16'h1623: data_out = 8'h39;
                    16'h1624: data_out = 8'h3A;
                    16'h1625: data_out = 8'h3B;
                    16'h1626: data_out = 8'h3C;
                    16'h1627: data_out = 8'h3D;
                    16'h1628: data_out = 8'h3E;
                    16'h1629: data_out = 8'h3F;
                    16'h162A: data_out = 8'h40;
                    16'h162B: data_out = 8'h41;
                    16'h162C: data_out = 8'h42;
                    16'h162D: data_out = 8'h43;
                    16'h162E: data_out = 8'h44;
                    16'h162F: data_out = 8'h45;
                    16'h1630: data_out = 8'h46;
                    16'h1631: data_out = 8'h47;
                    16'h1632: data_out = 8'h48;
                    16'h1633: data_out = 8'h49;
                    16'h1634: data_out = 8'h4A;
                    16'h1635: data_out = 8'h4B;
                    16'h1636: data_out = 8'h4C;
                    16'h1637: data_out = 8'h4D;
                    16'h1638: data_out = 8'h4E;
                    16'h1639: data_out = 8'h4F;
                    16'h163A: data_out = 8'h50;
                    16'h163B: data_out = 8'h51;
                    16'h163C: data_out = 8'h52;
                    16'h163D: data_out = 8'h53;
                    16'h163E: data_out = 8'h54;
                    16'h163F: data_out = 8'h55;
                    16'h1640: data_out = 8'h56;
                    16'h1641: data_out = 8'h57;
                    16'h1642: data_out = 8'h58;
                    16'h1643: data_out = 8'h59;
                    16'h1644: data_out = 8'h5A;
                    16'h1645: data_out = 8'h5B;
                    16'h1646: data_out = 8'h5C;
                    16'h1647: data_out = 8'h5D;
                    16'h1648: data_out = 8'h5E;
                    16'h1649: data_out = 8'h5F;
                    16'h164A: data_out = 8'h60;
                    16'h164B: data_out = 8'h61;
                    16'h164C: data_out = 8'h62;
                    16'h164D: data_out = 8'h63;
                    16'h164E: data_out = 8'h64;
                    16'h164F: data_out = 8'h65;
                    16'h1650: data_out = 8'h66;
                    16'h1651: data_out = 8'h67;
                    16'h1652: data_out = 8'h68;
                    16'h1653: data_out = 8'h69;
                    16'h1654: data_out = 8'h6A;
                    16'h1655: data_out = 8'h6B;
                    16'h1656: data_out = 8'h6C;
                    16'h1657: data_out = 8'h6D;
                    16'h1658: data_out = 8'h6E;
                    16'h1659: data_out = 8'h6F;
                    16'h165A: data_out = 8'h70;
                    16'h165B: data_out = 8'h71;
                    16'h165C: data_out = 8'h72;
                    16'h165D: data_out = 8'h73;
                    16'h165E: data_out = 8'h74;
                    16'h165F: data_out = 8'h75;
                    16'h1660: data_out = 8'h76;
                    16'h1661: data_out = 8'h77;
                    16'h1662: data_out = 8'h78;
                    16'h1663: data_out = 8'h79;
                    16'h1664: data_out = 8'h7A;
                    16'h1665: data_out = 8'h7B;
                    16'h1666: data_out = 8'h7C;
                    16'h1667: data_out = 8'h7D;
                    16'h1668: data_out = 8'h7E;
                    16'h1669: data_out = 8'h7F;
                    16'h166A: data_out = 8'h80;
                    16'h166B: data_out = 8'h81;
                    16'h166C: data_out = 8'h82;
                    16'h166D: data_out = 8'h83;
                    16'h166E: data_out = 8'h84;
                    16'h166F: data_out = 8'h85;
                    16'h1670: data_out = 8'h86;
                    16'h1671: data_out = 8'h87;
                    16'h1672: data_out = 8'h88;
                    16'h1673: data_out = 8'h89;
                    16'h1674: data_out = 8'h8A;
                    16'h1675: data_out = 8'h8B;
                    16'h1676: data_out = 8'h8C;
                    16'h1677: data_out = 8'h8D;
                    16'h1678: data_out = 8'h8E;
                    16'h1679: data_out = 8'h8F;
                    16'h167A: data_out = 8'h90;
                    16'h167B: data_out = 8'h91;
                    16'h167C: data_out = 8'h92;
                    16'h167D: data_out = 8'h93;
                    16'h167E: data_out = 8'h94;
                    16'h167F: data_out = 8'h95;
                    16'h1680: data_out = 8'h16;
                    16'h1681: data_out = 8'h15;
                    16'h1682: data_out = 8'h14;
                    16'h1683: data_out = 8'h13;
                    16'h1684: data_out = 8'h12;
                    16'h1685: data_out = 8'h11;
                    16'h1686: data_out = 8'h10;
                    16'h1687: data_out = 8'hF;
                    16'h1688: data_out = 8'hE;
                    16'h1689: data_out = 8'hD;
                    16'h168A: data_out = 8'hC;
                    16'h168B: data_out = 8'hB;
                    16'h168C: data_out = 8'hA;
                    16'h168D: data_out = 8'h9;
                    16'h168E: data_out = 8'h8;
                    16'h168F: data_out = 8'h7;
                    16'h1690: data_out = 8'h6;
                    16'h1691: data_out = 8'h5;
                    16'h1692: data_out = 8'h4;
                    16'h1693: data_out = 8'h3;
                    16'h1694: data_out = 8'h2;
                    16'h1695: data_out = 8'h1;
                    16'h1696: data_out = 8'h0;
                    16'h1697: data_out = 8'h81;
                    16'h1698: data_out = 8'h82;
                    16'h1699: data_out = 8'h83;
                    16'h169A: data_out = 8'h84;
                    16'h169B: data_out = 8'h85;
                    16'h169C: data_out = 8'h86;
                    16'h169D: data_out = 8'h87;
                    16'h169E: data_out = 8'h88;
                    16'h169F: data_out = 8'h89;
                    16'h16A0: data_out = 8'h8A;
                    16'h16A1: data_out = 8'h8B;
                    16'h16A2: data_out = 8'h8C;
                    16'h16A3: data_out = 8'h8D;
                    16'h16A4: data_out = 8'h8E;
                    16'h16A5: data_out = 8'h8F;
                    16'h16A6: data_out = 8'h90;
                    16'h16A7: data_out = 8'h91;
                    16'h16A8: data_out = 8'h92;
                    16'h16A9: data_out = 8'h93;
                    16'h16AA: data_out = 8'h94;
                    16'h16AB: data_out = 8'h95;
                    16'h16AC: data_out = 8'h96;
                    16'h16AD: data_out = 8'h97;
                    16'h16AE: data_out = 8'h98;
                    16'h16AF: data_out = 8'h99;
                    16'h16B0: data_out = 8'h9A;
                    16'h16B1: data_out = 8'h9B;
                    16'h16B2: data_out = 8'h9C;
                    16'h16B3: data_out = 8'h9D;
                    16'h16B4: data_out = 8'h9E;
                    16'h16B5: data_out = 8'h9F;
                    16'h16B6: data_out = 8'hA0;
                    16'h16B7: data_out = 8'hA1;
                    16'h16B8: data_out = 8'hA2;
                    16'h16B9: data_out = 8'hA3;
                    16'h16BA: data_out = 8'hA4;
                    16'h16BB: data_out = 8'hA5;
                    16'h16BC: data_out = 8'hA6;
                    16'h16BD: data_out = 8'hA7;
                    16'h16BE: data_out = 8'hA8;
                    16'h16BF: data_out = 8'hA9;
                    16'h16C0: data_out = 8'hAA;
                    16'h16C1: data_out = 8'hAB;
                    16'h16C2: data_out = 8'hAC;
                    16'h16C3: data_out = 8'hAD;
                    16'h16C4: data_out = 8'hAE;
                    16'h16C5: data_out = 8'hAF;
                    16'h16C6: data_out = 8'hB0;
                    16'h16C7: data_out = 8'hB1;
                    16'h16C8: data_out = 8'hB2;
                    16'h16C9: data_out = 8'hB3;
                    16'h16CA: data_out = 8'hB4;
                    16'h16CB: data_out = 8'hB5;
                    16'h16CC: data_out = 8'hB6;
                    16'h16CD: data_out = 8'hB7;
                    16'h16CE: data_out = 8'hB8;
                    16'h16CF: data_out = 8'hB9;
                    16'h16D0: data_out = 8'hBA;
                    16'h16D1: data_out = 8'hBB;
                    16'h16D2: data_out = 8'hBC;
                    16'h16D3: data_out = 8'hBD;
                    16'h16D4: data_out = 8'hBE;
                    16'h16D5: data_out = 8'hBF;
                    16'h16D6: data_out = 8'hC0;
                    16'h16D7: data_out = 8'hC1;
                    16'h16D8: data_out = 8'hC2;
                    16'h16D9: data_out = 8'hC3;
                    16'h16DA: data_out = 8'hC4;
                    16'h16DB: data_out = 8'hC5;
                    16'h16DC: data_out = 8'hC6;
                    16'h16DD: data_out = 8'hC7;
                    16'h16DE: data_out = 8'hC8;
                    16'h16DF: data_out = 8'hC9;
                    16'h16E0: data_out = 8'hCA;
                    16'h16E1: data_out = 8'hCB;
                    16'h16E2: data_out = 8'hCC;
                    16'h16E3: data_out = 8'hCD;
                    16'h16E4: data_out = 8'hCE;
                    16'h16E5: data_out = 8'hCF;
                    16'h16E6: data_out = 8'hD0;
                    16'h16E7: data_out = 8'hD1;
                    16'h16E8: data_out = 8'hD2;
                    16'h16E9: data_out = 8'hD3;
                    16'h16EA: data_out = 8'hD4;
                    16'h16EB: data_out = 8'hD5;
                    16'h16EC: data_out = 8'hD6;
                    16'h16ED: data_out = 8'hD7;
                    16'h16EE: data_out = 8'hD8;
                    16'h16EF: data_out = 8'hD9;
                    16'h16F0: data_out = 8'hDA;
                    16'h16F1: data_out = 8'hDB;
                    16'h16F2: data_out = 8'hDC;
                    16'h16F3: data_out = 8'hDD;
                    16'h16F4: data_out = 8'hDE;
                    16'h16F5: data_out = 8'hDF;
                    16'h16F6: data_out = 8'hE0;
                    16'h16F7: data_out = 8'hE1;
                    16'h16F8: data_out = 8'hE2;
                    16'h16F9: data_out = 8'hE3;
                    16'h16FA: data_out = 8'hE4;
                    16'h16FB: data_out = 8'hE5;
                    16'h16FC: data_out = 8'hE6;
                    16'h16FD: data_out = 8'hE7;
                    16'h16FE: data_out = 8'hE8;
                    16'h16FF: data_out = 8'hE9;
                    16'h1700: data_out = 8'h17;
                    16'h1701: data_out = 8'h18;
                    16'h1702: data_out = 8'h19;
                    16'h1703: data_out = 8'h1A;
                    16'h1704: data_out = 8'h1B;
                    16'h1705: data_out = 8'h1C;
                    16'h1706: data_out = 8'h1D;
                    16'h1707: data_out = 8'h1E;
                    16'h1708: data_out = 8'h1F;
                    16'h1709: data_out = 8'h20;
                    16'h170A: data_out = 8'h21;
                    16'h170B: data_out = 8'h22;
                    16'h170C: data_out = 8'h23;
                    16'h170D: data_out = 8'h24;
                    16'h170E: data_out = 8'h25;
                    16'h170F: data_out = 8'h26;
                    16'h1710: data_out = 8'h27;
                    16'h1711: data_out = 8'h28;
                    16'h1712: data_out = 8'h29;
                    16'h1713: data_out = 8'h2A;
                    16'h1714: data_out = 8'h2B;
                    16'h1715: data_out = 8'h2C;
                    16'h1716: data_out = 8'h2D;
                    16'h1717: data_out = 8'h2E;
                    16'h1718: data_out = 8'h2F;
                    16'h1719: data_out = 8'h30;
                    16'h171A: data_out = 8'h31;
                    16'h171B: data_out = 8'h32;
                    16'h171C: data_out = 8'h33;
                    16'h171D: data_out = 8'h34;
                    16'h171E: data_out = 8'h35;
                    16'h171F: data_out = 8'h36;
                    16'h1720: data_out = 8'h37;
                    16'h1721: data_out = 8'h38;
                    16'h1722: data_out = 8'h39;
                    16'h1723: data_out = 8'h3A;
                    16'h1724: data_out = 8'h3B;
                    16'h1725: data_out = 8'h3C;
                    16'h1726: data_out = 8'h3D;
                    16'h1727: data_out = 8'h3E;
                    16'h1728: data_out = 8'h3F;
                    16'h1729: data_out = 8'h40;
                    16'h172A: data_out = 8'h41;
                    16'h172B: data_out = 8'h42;
                    16'h172C: data_out = 8'h43;
                    16'h172D: data_out = 8'h44;
                    16'h172E: data_out = 8'h45;
                    16'h172F: data_out = 8'h46;
                    16'h1730: data_out = 8'h47;
                    16'h1731: data_out = 8'h48;
                    16'h1732: data_out = 8'h49;
                    16'h1733: data_out = 8'h4A;
                    16'h1734: data_out = 8'h4B;
                    16'h1735: data_out = 8'h4C;
                    16'h1736: data_out = 8'h4D;
                    16'h1737: data_out = 8'h4E;
                    16'h1738: data_out = 8'h4F;
                    16'h1739: data_out = 8'h50;
                    16'h173A: data_out = 8'h51;
                    16'h173B: data_out = 8'h52;
                    16'h173C: data_out = 8'h53;
                    16'h173D: data_out = 8'h54;
                    16'h173E: data_out = 8'h55;
                    16'h173F: data_out = 8'h56;
                    16'h1740: data_out = 8'h57;
                    16'h1741: data_out = 8'h58;
                    16'h1742: data_out = 8'h59;
                    16'h1743: data_out = 8'h5A;
                    16'h1744: data_out = 8'h5B;
                    16'h1745: data_out = 8'h5C;
                    16'h1746: data_out = 8'h5D;
                    16'h1747: data_out = 8'h5E;
                    16'h1748: data_out = 8'h5F;
                    16'h1749: data_out = 8'h60;
                    16'h174A: data_out = 8'h61;
                    16'h174B: data_out = 8'h62;
                    16'h174C: data_out = 8'h63;
                    16'h174D: data_out = 8'h64;
                    16'h174E: data_out = 8'h65;
                    16'h174F: data_out = 8'h66;
                    16'h1750: data_out = 8'h67;
                    16'h1751: data_out = 8'h68;
                    16'h1752: data_out = 8'h69;
                    16'h1753: data_out = 8'h6A;
                    16'h1754: data_out = 8'h6B;
                    16'h1755: data_out = 8'h6C;
                    16'h1756: data_out = 8'h6D;
                    16'h1757: data_out = 8'h6E;
                    16'h1758: data_out = 8'h6F;
                    16'h1759: data_out = 8'h70;
                    16'h175A: data_out = 8'h71;
                    16'h175B: data_out = 8'h72;
                    16'h175C: data_out = 8'h73;
                    16'h175D: data_out = 8'h74;
                    16'h175E: data_out = 8'h75;
                    16'h175F: data_out = 8'h76;
                    16'h1760: data_out = 8'h77;
                    16'h1761: data_out = 8'h78;
                    16'h1762: data_out = 8'h79;
                    16'h1763: data_out = 8'h7A;
                    16'h1764: data_out = 8'h7B;
                    16'h1765: data_out = 8'h7C;
                    16'h1766: data_out = 8'h7D;
                    16'h1767: data_out = 8'h7E;
                    16'h1768: data_out = 8'h7F;
                    16'h1769: data_out = 8'h80;
                    16'h176A: data_out = 8'h81;
                    16'h176B: data_out = 8'h82;
                    16'h176C: data_out = 8'h83;
                    16'h176D: data_out = 8'h84;
                    16'h176E: data_out = 8'h85;
                    16'h176F: data_out = 8'h86;
                    16'h1770: data_out = 8'h87;
                    16'h1771: data_out = 8'h88;
                    16'h1772: data_out = 8'h89;
                    16'h1773: data_out = 8'h8A;
                    16'h1774: data_out = 8'h8B;
                    16'h1775: data_out = 8'h8C;
                    16'h1776: data_out = 8'h8D;
                    16'h1777: data_out = 8'h8E;
                    16'h1778: data_out = 8'h8F;
                    16'h1779: data_out = 8'h90;
                    16'h177A: data_out = 8'h91;
                    16'h177B: data_out = 8'h92;
                    16'h177C: data_out = 8'h93;
                    16'h177D: data_out = 8'h94;
                    16'h177E: data_out = 8'h95;
                    16'h177F: data_out = 8'h96;
                    16'h1780: data_out = 8'h17;
                    16'h1781: data_out = 8'h16;
                    16'h1782: data_out = 8'h15;
                    16'h1783: data_out = 8'h14;
                    16'h1784: data_out = 8'h13;
                    16'h1785: data_out = 8'h12;
                    16'h1786: data_out = 8'h11;
                    16'h1787: data_out = 8'h10;
                    16'h1788: data_out = 8'hF;
                    16'h1789: data_out = 8'hE;
                    16'h178A: data_out = 8'hD;
                    16'h178B: data_out = 8'hC;
                    16'h178C: data_out = 8'hB;
                    16'h178D: data_out = 8'hA;
                    16'h178E: data_out = 8'h9;
                    16'h178F: data_out = 8'h8;
                    16'h1790: data_out = 8'h7;
                    16'h1791: data_out = 8'h6;
                    16'h1792: data_out = 8'h5;
                    16'h1793: data_out = 8'h4;
                    16'h1794: data_out = 8'h3;
                    16'h1795: data_out = 8'h2;
                    16'h1796: data_out = 8'h1;
                    16'h1797: data_out = 8'h0;
                    16'h1798: data_out = 8'h81;
                    16'h1799: data_out = 8'h82;
                    16'h179A: data_out = 8'h83;
                    16'h179B: data_out = 8'h84;
                    16'h179C: data_out = 8'h85;
                    16'h179D: data_out = 8'h86;
                    16'h179E: data_out = 8'h87;
                    16'h179F: data_out = 8'h88;
                    16'h17A0: data_out = 8'h89;
                    16'h17A1: data_out = 8'h8A;
                    16'h17A2: data_out = 8'h8B;
                    16'h17A3: data_out = 8'h8C;
                    16'h17A4: data_out = 8'h8D;
                    16'h17A5: data_out = 8'h8E;
                    16'h17A6: data_out = 8'h8F;
                    16'h17A7: data_out = 8'h90;
                    16'h17A8: data_out = 8'h91;
                    16'h17A9: data_out = 8'h92;
                    16'h17AA: data_out = 8'h93;
                    16'h17AB: data_out = 8'h94;
                    16'h17AC: data_out = 8'h95;
                    16'h17AD: data_out = 8'h96;
                    16'h17AE: data_out = 8'h97;
                    16'h17AF: data_out = 8'h98;
                    16'h17B0: data_out = 8'h99;
                    16'h17B1: data_out = 8'h9A;
                    16'h17B2: data_out = 8'h9B;
                    16'h17B3: data_out = 8'h9C;
                    16'h17B4: data_out = 8'h9D;
                    16'h17B5: data_out = 8'h9E;
                    16'h17B6: data_out = 8'h9F;
                    16'h17B7: data_out = 8'hA0;
                    16'h17B8: data_out = 8'hA1;
                    16'h17B9: data_out = 8'hA2;
                    16'h17BA: data_out = 8'hA3;
                    16'h17BB: data_out = 8'hA4;
                    16'h17BC: data_out = 8'hA5;
                    16'h17BD: data_out = 8'hA6;
                    16'h17BE: data_out = 8'hA7;
                    16'h17BF: data_out = 8'hA8;
                    16'h17C0: data_out = 8'hA9;
                    16'h17C1: data_out = 8'hAA;
                    16'h17C2: data_out = 8'hAB;
                    16'h17C3: data_out = 8'hAC;
                    16'h17C4: data_out = 8'hAD;
                    16'h17C5: data_out = 8'hAE;
                    16'h17C6: data_out = 8'hAF;
                    16'h17C7: data_out = 8'hB0;
                    16'h17C8: data_out = 8'hB1;
                    16'h17C9: data_out = 8'hB2;
                    16'h17CA: data_out = 8'hB3;
                    16'h17CB: data_out = 8'hB4;
                    16'h17CC: data_out = 8'hB5;
                    16'h17CD: data_out = 8'hB6;
                    16'h17CE: data_out = 8'hB7;
                    16'h17CF: data_out = 8'hB8;
                    16'h17D0: data_out = 8'hB9;
                    16'h17D1: data_out = 8'hBA;
                    16'h17D2: data_out = 8'hBB;
                    16'h17D3: data_out = 8'hBC;
                    16'h17D4: data_out = 8'hBD;
                    16'h17D5: data_out = 8'hBE;
                    16'h17D6: data_out = 8'hBF;
                    16'h17D7: data_out = 8'hC0;
                    16'h17D8: data_out = 8'hC1;
                    16'h17D9: data_out = 8'hC2;
                    16'h17DA: data_out = 8'hC3;
                    16'h17DB: data_out = 8'hC4;
                    16'h17DC: data_out = 8'hC5;
                    16'h17DD: data_out = 8'hC6;
                    16'h17DE: data_out = 8'hC7;
                    16'h17DF: data_out = 8'hC8;
                    16'h17E0: data_out = 8'hC9;
                    16'h17E1: data_out = 8'hCA;
                    16'h17E2: data_out = 8'hCB;
                    16'h17E3: data_out = 8'hCC;
                    16'h17E4: data_out = 8'hCD;
                    16'h17E5: data_out = 8'hCE;
                    16'h17E6: data_out = 8'hCF;
                    16'h17E7: data_out = 8'hD0;
                    16'h17E8: data_out = 8'hD1;
                    16'h17E9: data_out = 8'hD2;
                    16'h17EA: data_out = 8'hD3;
                    16'h17EB: data_out = 8'hD4;
                    16'h17EC: data_out = 8'hD5;
                    16'h17ED: data_out = 8'hD6;
                    16'h17EE: data_out = 8'hD7;
                    16'h17EF: data_out = 8'hD8;
                    16'h17F0: data_out = 8'hD9;
                    16'h17F1: data_out = 8'hDA;
                    16'h17F2: data_out = 8'hDB;
                    16'h17F3: data_out = 8'hDC;
                    16'h17F4: data_out = 8'hDD;
                    16'h17F5: data_out = 8'hDE;
                    16'h17F6: data_out = 8'hDF;
                    16'h17F7: data_out = 8'hE0;
                    16'h17F8: data_out = 8'hE1;
                    16'h17F9: data_out = 8'hE2;
                    16'h17FA: data_out = 8'hE3;
                    16'h17FB: data_out = 8'hE4;
                    16'h17FC: data_out = 8'hE5;
                    16'h17FD: data_out = 8'hE6;
                    16'h17FE: data_out = 8'hE7;
                    16'h17FF: data_out = 8'hE8;
                    16'h1800: data_out = 8'h18;
                    16'h1801: data_out = 8'h19;
                    16'h1802: data_out = 8'h1A;
                    16'h1803: data_out = 8'h1B;
                    16'h1804: data_out = 8'h1C;
                    16'h1805: data_out = 8'h1D;
                    16'h1806: data_out = 8'h1E;
                    16'h1807: data_out = 8'h1F;
                    16'h1808: data_out = 8'h20;
                    16'h1809: data_out = 8'h21;
                    16'h180A: data_out = 8'h22;
                    16'h180B: data_out = 8'h23;
                    16'h180C: data_out = 8'h24;
                    16'h180D: data_out = 8'h25;
                    16'h180E: data_out = 8'h26;
                    16'h180F: data_out = 8'h27;
                    16'h1810: data_out = 8'h28;
                    16'h1811: data_out = 8'h29;
                    16'h1812: data_out = 8'h2A;
                    16'h1813: data_out = 8'h2B;
                    16'h1814: data_out = 8'h2C;
                    16'h1815: data_out = 8'h2D;
                    16'h1816: data_out = 8'h2E;
                    16'h1817: data_out = 8'h2F;
                    16'h1818: data_out = 8'h30;
                    16'h1819: data_out = 8'h31;
                    16'h181A: data_out = 8'h32;
                    16'h181B: data_out = 8'h33;
                    16'h181C: data_out = 8'h34;
                    16'h181D: data_out = 8'h35;
                    16'h181E: data_out = 8'h36;
                    16'h181F: data_out = 8'h37;
                    16'h1820: data_out = 8'h38;
                    16'h1821: data_out = 8'h39;
                    16'h1822: data_out = 8'h3A;
                    16'h1823: data_out = 8'h3B;
                    16'h1824: data_out = 8'h3C;
                    16'h1825: data_out = 8'h3D;
                    16'h1826: data_out = 8'h3E;
                    16'h1827: data_out = 8'h3F;
                    16'h1828: data_out = 8'h40;
                    16'h1829: data_out = 8'h41;
                    16'h182A: data_out = 8'h42;
                    16'h182B: data_out = 8'h43;
                    16'h182C: data_out = 8'h44;
                    16'h182D: data_out = 8'h45;
                    16'h182E: data_out = 8'h46;
                    16'h182F: data_out = 8'h47;
                    16'h1830: data_out = 8'h48;
                    16'h1831: data_out = 8'h49;
                    16'h1832: data_out = 8'h4A;
                    16'h1833: data_out = 8'h4B;
                    16'h1834: data_out = 8'h4C;
                    16'h1835: data_out = 8'h4D;
                    16'h1836: data_out = 8'h4E;
                    16'h1837: data_out = 8'h4F;
                    16'h1838: data_out = 8'h50;
                    16'h1839: data_out = 8'h51;
                    16'h183A: data_out = 8'h52;
                    16'h183B: data_out = 8'h53;
                    16'h183C: data_out = 8'h54;
                    16'h183D: data_out = 8'h55;
                    16'h183E: data_out = 8'h56;
                    16'h183F: data_out = 8'h57;
                    16'h1840: data_out = 8'h58;
                    16'h1841: data_out = 8'h59;
                    16'h1842: data_out = 8'h5A;
                    16'h1843: data_out = 8'h5B;
                    16'h1844: data_out = 8'h5C;
                    16'h1845: data_out = 8'h5D;
                    16'h1846: data_out = 8'h5E;
                    16'h1847: data_out = 8'h5F;
                    16'h1848: data_out = 8'h60;
                    16'h1849: data_out = 8'h61;
                    16'h184A: data_out = 8'h62;
                    16'h184B: data_out = 8'h63;
                    16'h184C: data_out = 8'h64;
                    16'h184D: data_out = 8'h65;
                    16'h184E: data_out = 8'h66;
                    16'h184F: data_out = 8'h67;
                    16'h1850: data_out = 8'h68;
                    16'h1851: data_out = 8'h69;
                    16'h1852: data_out = 8'h6A;
                    16'h1853: data_out = 8'h6B;
                    16'h1854: data_out = 8'h6C;
                    16'h1855: data_out = 8'h6D;
                    16'h1856: data_out = 8'h6E;
                    16'h1857: data_out = 8'h6F;
                    16'h1858: data_out = 8'h70;
                    16'h1859: data_out = 8'h71;
                    16'h185A: data_out = 8'h72;
                    16'h185B: data_out = 8'h73;
                    16'h185C: data_out = 8'h74;
                    16'h185D: data_out = 8'h75;
                    16'h185E: data_out = 8'h76;
                    16'h185F: data_out = 8'h77;
                    16'h1860: data_out = 8'h78;
                    16'h1861: data_out = 8'h79;
                    16'h1862: data_out = 8'h7A;
                    16'h1863: data_out = 8'h7B;
                    16'h1864: data_out = 8'h7C;
                    16'h1865: data_out = 8'h7D;
                    16'h1866: data_out = 8'h7E;
                    16'h1867: data_out = 8'h7F;
                    16'h1868: data_out = 8'h80;
                    16'h1869: data_out = 8'h81;
                    16'h186A: data_out = 8'h82;
                    16'h186B: data_out = 8'h83;
                    16'h186C: data_out = 8'h84;
                    16'h186D: data_out = 8'h85;
                    16'h186E: data_out = 8'h86;
                    16'h186F: data_out = 8'h87;
                    16'h1870: data_out = 8'h88;
                    16'h1871: data_out = 8'h89;
                    16'h1872: data_out = 8'h8A;
                    16'h1873: data_out = 8'h8B;
                    16'h1874: data_out = 8'h8C;
                    16'h1875: data_out = 8'h8D;
                    16'h1876: data_out = 8'h8E;
                    16'h1877: data_out = 8'h8F;
                    16'h1878: data_out = 8'h90;
                    16'h1879: data_out = 8'h91;
                    16'h187A: data_out = 8'h92;
                    16'h187B: data_out = 8'h93;
                    16'h187C: data_out = 8'h94;
                    16'h187D: data_out = 8'h95;
                    16'h187E: data_out = 8'h96;
                    16'h187F: data_out = 8'h97;
                    16'h1880: data_out = 8'h18;
                    16'h1881: data_out = 8'h17;
                    16'h1882: data_out = 8'h16;
                    16'h1883: data_out = 8'h15;
                    16'h1884: data_out = 8'h14;
                    16'h1885: data_out = 8'h13;
                    16'h1886: data_out = 8'h12;
                    16'h1887: data_out = 8'h11;
                    16'h1888: data_out = 8'h10;
                    16'h1889: data_out = 8'hF;
                    16'h188A: data_out = 8'hE;
                    16'h188B: data_out = 8'hD;
                    16'h188C: data_out = 8'hC;
                    16'h188D: data_out = 8'hB;
                    16'h188E: data_out = 8'hA;
                    16'h188F: data_out = 8'h9;
                    16'h1890: data_out = 8'h8;
                    16'h1891: data_out = 8'h7;
                    16'h1892: data_out = 8'h6;
                    16'h1893: data_out = 8'h5;
                    16'h1894: data_out = 8'h4;
                    16'h1895: data_out = 8'h3;
                    16'h1896: data_out = 8'h2;
                    16'h1897: data_out = 8'h1;
                    16'h1898: data_out = 8'h0;
                    16'h1899: data_out = 8'h81;
                    16'h189A: data_out = 8'h82;
                    16'h189B: data_out = 8'h83;
                    16'h189C: data_out = 8'h84;
                    16'h189D: data_out = 8'h85;
                    16'h189E: data_out = 8'h86;
                    16'h189F: data_out = 8'h87;
                    16'h18A0: data_out = 8'h88;
                    16'h18A1: data_out = 8'h89;
                    16'h18A2: data_out = 8'h8A;
                    16'h18A3: data_out = 8'h8B;
                    16'h18A4: data_out = 8'h8C;
                    16'h18A5: data_out = 8'h8D;
                    16'h18A6: data_out = 8'h8E;
                    16'h18A7: data_out = 8'h8F;
                    16'h18A8: data_out = 8'h90;
                    16'h18A9: data_out = 8'h91;
                    16'h18AA: data_out = 8'h92;
                    16'h18AB: data_out = 8'h93;
                    16'h18AC: data_out = 8'h94;
                    16'h18AD: data_out = 8'h95;
                    16'h18AE: data_out = 8'h96;
                    16'h18AF: data_out = 8'h97;
                    16'h18B0: data_out = 8'h98;
                    16'h18B1: data_out = 8'h99;
                    16'h18B2: data_out = 8'h9A;
                    16'h18B3: data_out = 8'h9B;
                    16'h18B4: data_out = 8'h9C;
                    16'h18B5: data_out = 8'h9D;
                    16'h18B6: data_out = 8'h9E;
                    16'h18B7: data_out = 8'h9F;
                    16'h18B8: data_out = 8'hA0;
                    16'h18B9: data_out = 8'hA1;
                    16'h18BA: data_out = 8'hA2;
                    16'h18BB: data_out = 8'hA3;
                    16'h18BC: data_out = 8'hA4;
                    16'h18BD: data_out = 8'hA5;
                    16'h18BE: data_out = 8'hA6;
                    16'h18BF: data_out = 8'hA7;
                    16'h18C0: data_out = 8'hA8;
                    16'h18C1: data_out = 8'hA9;
                    16'h18C2: data_out = 8'hAA;
                    16'h18C3: data_out = 8'hAB;
                    16'h18C4: data_out = 8'hAC;
                    16'h18C5: data_out = 8'hAD;
                    16'h18C6: data_out = 8'hAE;
                    16'h18C7: data_out = 8'hAF;
                    16'h18C8: data_out = 8'hB0;
                    16'h18C9: data_out = 8'hB1;
                    16'h18CA: data_out = 8'hB2;
                    16'h18CB: data_out = 8'hB3;
                    16'h18CC: data_out = 8'hB4;
                    16'h18CD: data_out = 8'hB5;
                    16'h18CE: data_out = 8'hB6;
                    16'h18CF: data_out = 8'hB7;
                    16'h18D0: data_out = 8'hB8;
                    16'h18D1: data_out = 8'hB9;
                    16'h18D2: data_out = 8'hBA;
                    16'h18D3: data_out = 8'hBB;
                    16'h18D4: data_out = 8'hBC;
                    16'h18D5: data_out = 8'hBD;
                    16'h18D6: data_out = 8'hBE;
                    16'h18D7: data_out = 8'hBF;
                    16'h18D8: data_out = 8'hC0;
                    16'h18D9: data_out = 8'hC1;
                    16'h18DA: data_out = 8'hC2;
                    16'h18DB: data_out = 8'hC3;
                    16'h18DC: data_out = 8'hC4;
                    16'h18DD: data_out = 8'hC5;
                    16'h18DE: data_out = 8'hC6;
                    16'h18DF: data_out = 8'hC7;
                    16'h18E0: data_out = 8'hC8;
                    16'h18E1: data_out = 8'hC9;
                    16'h18E2: data_out = 8'hCA;
                    16'h18E3: data_out = 8'hCB;
                    16'h18E4: data_out = 8'hCC;
                    16'h18E5: data_out = 8'hCD;
                    16'h18E6: data_out = 8'hCE;
                    16'h18E7: data_out = 8'hCF;
                    16'h18E8: data_out = 8'hD0;
                    16'h18E9: data_out = 8'hD1;
                    16'h18EA: data_out = 8'hD2;
                    16'h18EB: data_out = 8'hD3;
                    16'h18EC: data_out = 8'hD4;
                    16'h18ED: data_out = 8'hD5;
                    16'h18EE: data_out = 8'hD6;
                    16'h18EF: data_out = 8'hD7;
                    16'h18F0: data_out = 8'hD8;
                    16'h18F1: data_out = 8'hD9;
                    16'h18F2: data_out = 8'hDA;
                    16'h18F3: data_out = 8'hDB;
                    16'h18F4: data_out = 8'hDC;
                    16'h18F5: data_out = 8'hDD;
                    16'h18F6: data_out = 8'hDE;
                    16'h18F7: data_out = 8'hDF;
                    16'h18F8: data_out = 8'hE0;
                    16'h18F9: data_out = 8'hE1;
                    16'h18FA: data_out = 8'hE2;
                    16'h18FB: data_out = 8'hE3;
                    16'h18FC: data_out = 8'hE4;
                    16'h18FD: data_out = 8'hE5;
                    16'h18FE: data_out = 8'hE6;
                    16'h18FF: data_out = 8'hE7;
                    16'h1900: data_out = 8'h19;
                    16'h1901: data_out = 8'h1A;
                    16'h1902: data_out = 8'h1B;
                    16'h1903: data_out = 8'h1C;
                    16'h1904: data_out = 8'h1D;
                    16'h1905: data_out = 8'h1E;
                    16'h1906: data_out = 8'h1F;
                    16'h1907: data_out = 8'h20;
                    16'h1908: data_out = 8'h21;
                    16'h1909: data_out = 8'h22;
                    16'h190A: data_out = 8'h23;
                    16'h190B: data_out = 8'h24;
                    16'h190C: data_out = 8'h25;
                    16'h190D: data_out = 8'h26;
                    16'h190E: data_out = 8'h27;
                    16'h190F: data_out = 8'h28;
                    16'h1910: data_out = 8'h29;
                    16'h1911: data_out = 8'h2A;
                    16'h1912: data_out = 8'h2B;
                    16'h1913: data_out = 8'h2C;
                    16'h1914: data_out = 8'h2D;
                    16'h1915: data_out = 8'h2E;
                    16'h1916: data_out = 8'h2F;
                    16'h1917: data_out = 8'h30;
                    16'h1918: data_out = 8'h31;
                    16'h1919: data_out = 8'h32;
                    16'h191A: data_out = 8'h33;
                    16'h191B: data_out = 8'h34;
                    16'h191C: data_out = 8'h35;
                    16'h191D: data_out = 8'h36;
                    16'h191E: data_out = 8'h37;
                    16'h191F: data_out = 8'h38;
                    16'h1920: data_out = 8'h39;
                    16'h1921: data_out = 8'h3A;
                    16'h1922: data_out = 8'h3B;
                    16'h1923: data_out = 8'h3C;
                    16'h1924: data_out = 8'h3D;
                    16'h1925: data_out = 8'h3E;
                    16'h1926: data_out = 8'h3F;
                    16'h1927: data_out = 8'h40;
                    16'h1928: data_out = 8'h41;
                    16'h1929: data_out = 8'h42;
                    16'h192A: data_out = 8'h43;
                    16'h192B: data_out = 8'h44;
                    16'h192C: data_out = 8'h45;
                    16'h192D: data_out = 8'h46;
                    16'h192E: data_out = 8'h47;
                    16'h192F: data_out = 8'h48;
                    16'h1930: data_out = 8'h49;
                    16'h1931: data_out = 8'h4A;
                    16'h1932: data_out = 8'h4B;
                    16'h1933: data_out = 8'h4C;
                    16'h1934: data_out = 8'h4D;
                    16'h1935: data_out = 8'h4E;
                    16'h1936: data_out = 8'h4F;
                    16'h1937: data_out = 8'h50;
                    16'h1938: data_out = 8'h51;
                    16'h1939: data_out = 8'h52;
                    16'h193A: data_out = 8'h53;
                    16'h193B: data_out = 8'h54;
                    16'h193C: data_out = 8'h55;
                    16'h193D: data_out = 8'h56;
                    16'h193E: data_out = 8'h57;
                    16'h193F: data_out = 8'h58;
                    16'h1940: data_out = 8'h59;
                    16'h1941: data_out = 8'h5A;
                    16'h1942: data_out = 8'h5B;
                    16'h1943: data_out = 8'h5C;
                    16'h1944: data_out = 8'h5D;
                    16'h1945: data_out = 8'h5E;
                    16'h1946: data_out = 8'h5F;
                    16'h1947: data_out = 8'h60;
                    16'h1948: data_out = 8'h61;
                    16'h1949: data_out = 8'h62;
                    16'h194A: data_out = 8'h63;
                    16'h194B: data_out = 8'h64;
                    16'h194C: data_out = 8'h65;
                    16'h194D: data_out = 8'h66;
                    16'h194E: data_out = 8'h67;
                    16'h194F: data_out = 8'h68;
                    16'h1950: data_out = 8'h69;
                    16'h1951: data_out = 8'h6A;
                    16'h1952: data_out = 8'h6B;
                    16'h1953: data_out = 8'h6C;
                    16'h1954: data_out = 8'h6D;
                    16'h1955: data_out = 8'h6E;
                    16'h1956: data_out = 8'h6F;
                    16'h1957: data_out = 8'h70;
                    16'h1958: data_out = 8'h71;
                    16'h1959: data_out = 8'h72;
                    16'h195A: data_out = 8'h73;
                    16'h195B: data_out = 8'h74;
                    16'h195C: data_out = 8'h75;
                    16'h195D: data_out = 8'h76;
                    16'h195E: data_out = 8'h77;
                    16'h195F: data_out = 8'h78;
                    16'h1960: data_out = 8'h79;
                    16'h1961: data_out = 8'h7A;
                    16'h1962: data_out = 8'h7B;
                    16'h1963: data_out = 8'h7C;
                    16'h1964: data_out = 8'h7D;
                    16'h1965: data_out = 8'h7E;
                    16'h1966: data_out = 8'h7F;
                    16'h1967: data_out = 8'h80;
                    16'h1968: data_out = 8'h81;
                    16'h1969: data_out = 8'h82;
                    16'h196A: data_out = 8'h83;
                    16'h196B: data_out = 8'h84;
                    16'h196C: data_out = 8'h85;
                    16'h196D: data_out = 8'h86;
                    16'h196E: data_out = 8'h87;
                    16'h196F: data_out = 8'h88;
                    16'h1970: data_out = 8'h89;
                    16'h1971: data_out = 8'h8A;
                    16'h1972: data_out = 8'h8B;
                    16'h1973: data_out = 8'h8C;
                    16'h1974: data_out = 8'h8D;
                    16'h1975: data_out = 8'h8E;
                    16'h1976: data_out = 8'h8F;
                    16'h1977: data_out = 8'h90;
                    16'h1978: data_out = 8'h91;
                    16'h1979: data_out = 8'h92;
                    16'h197A: data_out = 8'h93;
                    16'h197B: data_out = 8'h94;
                    16'h197C: data_out = 8'h95;
                    16'h197D: data_out = 8'h96;
                    16'h197E: data_out = 8'h97;
                    16'h197F: data_out = 8'h98;
                    16'h1980: data_out = 8'h19;
                    16'h1981: data_out = 8'h18;
                    16'h1982: data_out = 8'h17;
                    16'h1983: data_out = 8'h16;
                    16'h1984: data_out = 8'h15;
                    16'h1985: data_out = 8'h14;
                    16'h1986: data_out = 8'h13;
                    16'h1987: data_out = 8'h12;
                    16'h1988: data_out = 8'h11;
                    16'h1989: data_out = 8'h10;
                    16'h198A: data_out = 8'hF;
                    16'h198B: data_out = 8'hE;
                    16'h198C: data_out = 8'hD;
                    16'h198D: data_out = 8'hC;
                    16'h198E: data_out = 8'hB;
                    16'h198F: data_out = 8'hA;
                    16'h1990: data_out = 8'h9;
                    16'h1991: data_out = 8'h8;
                    16'h1992: data_out = 8'h7;
                    16'h1993: data_out = 8'h6;
                    16'h1994: data_out = 8'h5;
                    16'h1995: data_out = 8'h4;
                    16'h1996: data_out = 8'h3;
                    16'h1997: data_out = 8'h2;
                    16'h1998: data_out = 8'h1;
                    16'h1999: data_out = 8'h0;
                    16'h199A: data_out = 8'h81;
                    16'h199B: data_out = 8'h82;
                    16'h199C: data_out = 8'h83;
                    16'h199D: data_out = 8'h84;
                    16'h199E: data_out = 8'h85;
                    16'h199F: data_out = 8'h86;
                    16'h19A0: data_out = 8'h87;
                    16'h19A1: data_out = 8'h88;
                    16'h19A2: data_out = 8'h89;
                    16'h19A3: data_out = 8'h8A;
                    16'h19A4: data_out = 8'h8B;
                    16'h19A5: data_out = 8'h8C;
                    16'h19A6: data_out = 8'h8D;
                    16'h19A7: data_out = 8'h8E;
                    16'h19A8: data_out = 8'h8F;
                    16'h19A9: data_out = 8'h90;
                    16'h19AA: data_out = 8'h91;
                    16'h19AB: data_out = 8'h92;
                    16'h19AC: data_out = 8'h93;
                    16'h19AD: data_out = 8'h94;
                    16'h19AE: data_out = 8'h95;
                    16'h19AF: data_out = 8'h96;
                    16'h19B0: data_out = 8'h97;
                    16'h19B1: data_out = 8'h98;
                    16'h19B2: data_out = 8'h99;
                    16'h19B3: data_out = 8'h9A;
                    16'h19B4: data_out = 8'h9B;
                    16'h19B5: data_out = 8'h9C;
                    16'h19B6: data_out = 8'h9D;
                    16'h19B7: data_out = 8'h9E;
                    16'h19B8: data_out = 8'h9F;
                    16'h19B9: data_out = 8'hA0;
                    16'h19BA: data_out = 8'hA1;
                    16'h19BB: data_out = 8'hA2;
                    16'h19BC: data_out = 8'hA3;
                    16'h19BD: data_out = 8'hA4;
                    16'h19BE: data_out = 8'hA5;
                    16'h19BF: data_out = 8'hA6;
                    16'h19C0: data_out = 8'hA7;
                    16'h19C1: data_out = 8'hA8;
                    16'h19C2: data_out = 8'hA9;
                    16'h19C3: data_out = 8'hAA;
                    16'h19C4: data_out = 8'hAB;
                    16'h19C5: data_out = 8'hAC;
                    16'h19C6: data_out = 8'hAD;
                    16'h19C7: data_out = 8'hAE;
                    16'h19C8: data_out = 8'hAF;
                    16'h19C9: data_out = 8'hB0;
                    16'h19CA: data_out = 8'hB1;
                    16'h19CB: data_out = 8'hB2;
                    16'h19CC: data_out = 8'hB3;
                    16'h19CD: data_out = 8'hB4;
                    16'h19CE: data_out = 8'hB5;
                    16'h19CF: data_out = 8'hB6;
                    16'h19D0: data_out = 8'hB7;
                    16'h19D1: data_out = 8'hB8;
                    16'h19D2: data_out = 8'hB9;
                    16'h19D3: data_out = 8'hBA;
                    16'h19D4: data_out = 8'hBB;
                    16'h19D5: data_out = 8'hBC;
                    16'h19D6: data_out = 8'hBD;
                    16'h19D7: data_out = 8'hBE;
                    16'h19D8: data_out = 8'hBF;
                    16'h19D9: data_out = 8'hC0;
                    16'h19DA: data_out = 8'hC1;
                    16'h19DB: data_out = 8'hC2;
                    16'h19DC: data_out = 8'hC3;
                    16'h19DD: data_out = 8'hC4;
                    16'h19DE: data_out = 8'hC5;
                    16'h19DF: data_out = 8'hC6;
                    16'h19E0: data_out = 8'hC7;
                    16'h19E1: data_out = 8'hC8;
                    16'h19E2: data_out = 8'hC9;
                    16'h19E3: data_out = 8'hCA;
                    16'h19E4: data_out = 8'hCB;
                    16'h19E5: data_out = 8'hCC;
                    16'h19E6: data_out = 8'hCD;
                    16'h19E7: data_out = 8'hCE;
                    16'h19E8: data_out = 8'hCF;
                    16'h19E9: data_out = 8'hD0;
                    16'h19EA: data_out = 8'hD1;
                    16'h19EB: data_out = 8'hD2;
                    16'h19EC: data_out = 8'hD3;
                    16'h19ED: data_out = 8'hD4;
                    16'h19EE: data_out = 8'hD5;
                    16'h19EF: data_out = 8'hD6;
                    16'h19F0: data_out = 8'hD7;
                    16'h19F1: data_out = 8'hD8;
                    16'h19F2: data_out = 8'hD9;
                    16'h19F3: data_out = 8'hDA;
                    16'h19F4: data_out = 8'hDB;
                    16'h19F5: data_out = 8'hDC;
                    16'h19F6: data_out = 8'hDD;
                    16'h19F7: data_out = 8'hDE;
                    16'h19F8: data_out = 8'hDF;
                    16'h19F9: data_out = 8'hE0;
                    16'h19FA: data_out = 8'hE1;
                    16'h19FB: data_out = 8'hE2;
                    16'h19FC: data_out = 8'hE3;
                    16'h19FD: data_out = 8'hE4;
                    16'h19FE: data_out = 8'hE5;
                    16'h19FF: data_out = 8'hE6;
                    16'h1A00: data_out = 8'h1A;
                    16'h1A01: data_out = 8'h1B;
                    16'h1A02: data_out = 8'h1C;
                    16'h1A03: data_out = 8'h1D;
                    16'h1A04: data_out = 8'h1E;
                    16'h1A05: data_out = 8'h1F;
                    16'h1A06: data_out = 8'h20;
                    16'h1A07: data_out = 8'h21;
                    16'h1A08: data_out = 8'h22;
                    16'h1A09: data_out = 8'h23;
                    16'h1A0A: data_out = 8'h24;
                    16'h1A0B: data_out = 8'h25;
                    16'h1A0C: data_out = 8'h26;
                    16'h1A0D: data_out = 8'h27;
                    16'h1A0E: data_out = 8'h28;
                    16'h1A0F: data_out = 8'h29;
                    16'h1A10: data_out = 8'h2A;
                    16'h1A11: data_out = 8'h2B;
                    16'h1A12: data_out = 8'h2C;
                    16'h1A13: data_out = 8'h2D;
                    16'h1A14: data_out = 8'h2E;
                    16'h1A15: data_out = 8'h2F;
                    16'h1A16: data_out = 8'h30;
                    16'h1A17: data_out = 8'h31;
                    16'h1A18: data_out = 8'h32;
                    16'h1A19: data_out = 8'h33;
                    16'h1A1A: data_out = 8'h34;
                    16'h1A1B: data_out = 8'h35;
                    16'h1A1C: data_out = 8'h36;
                    16'h1A1D: data_out = 8'h37;
                    16'h1A1E: data_out = 8'h38;
                    16'h1A1F: data_out = 8'h39;
                    16'h1A20: data_out = 8'h3A;
                    16'h1A21: data_out = 8'h3B;
                    16'h1A22: data_out = 8'h3C;
                    16'h1A23: data_out = 8'h3D;
                    16'h1A24: data_out = 8'h3E;
                    16'h1A25: data_out = 8'h3F;
                    16'h1A26: data_out = 8'h40;
                    16'h1A27: data_out = 8'h41;
                    16'h1A28: data_out = 8'h42;
                    16'h1A29: data_out = 8'h43;
                    16'h1A2A: data_out = 8'h44;
                    16'h1A2B: data_out = 8'h45;
                    16'h1A2C: data_out = 8'h46;
                    16'h1A2D: data_out = 8'h47;
                    16'h1A2E: data_out = 8'h48;
                    16'h1A2F: data_out = 8'h49;
                    16'h1A30: data_out = 8'h4A;
                    16'h1A31: data_out = 8'h4B;
                    16'h1A32: data_out = 8'h4C;
                    16'h1A33: data_out = 8'h4D;
                    16'h1A34: data_out = 8'h4E;
                    16'h1A35: data_out = 8'h4F;
                    16'h1A36: data_out = 8'h50;
                    16'h1A37: data_out = 8'h51;
                    16'h1A38: data_out = 8'h52;
                    16'h1A39: data_out = 8'h53;
                    16'h1A3A: data_out = 8'h54;
                    16'h1A3B: data_out = 8'h55;
                    16'h1A3C: data_out = 8'h56;
                    16'h1A3D: data_out = 8'h57;
                    16'h1A3E: data_out = 8'h58;
                    16'h1A3F: data_out = 8'h59;
                    16'h1A40: data_out = 8'h5A;
                    16'h1A41: data_out = 8'h5B;
                    16'h1A42: data_out = 8'h5C;
                    16'h1A43: data_out = 8'h5D;
                    16'h1A44: data_out = 8'h5E;
                    16'h1A45: data_out = 8'h5F;
                    16'h1A46: data_out = 8'h60;
                    16'h1A47: data_out = 8'h61;
                    16'h1A48: data_out = 8'h62;
                    16'h1A49: data_out = 8'h63;
                    16'h1A4A: data_out = 8'h64;
                    16'h1A4B: data_out = 8'h65;
                    16'h1A4C: data_out = 8'h66;
                    16'h1A4D: data_out = 8'h67;
                    16'h1A4E: data_out = 8'h68;
                    16'h1A4F: data_out = 8'h69;
                    16'h1A50: data_out = 8'h6A;
                    16'h1A51: data_out = 8'h6B;
                    16'h1A52: data_out = 8'h6C;
                    16'h1A53: data_out = 8'h6D;
                    16'h1A54: data_out = 8'h6E;
                    16'h1A55: data_out = 8'h6F;
                    16'h1A56: data_out = 8'h70;
                    16'h1A57: data_out = 8'h71;
                    16'h1A58: data_out = 8'h72;
                    16'h1A59: data_out = 8'h73;
                    16'h1A5A: data_out = 8'h74;
                    16'h1A5B: data_out = 8'h75;
                    16'h1A5C: data_out = 8'h76;
                    16'h1A5D: data_out = 8'h77;
                    16'h1A5E: data_out = 8'h78;
                    16'h1A5F: data_out = 8'h79;
                    16'h1A60: data_out = 8'h7A;
                    16'h1A61: data_out = 8'h7B;
                    16'h1A62: data_out = 8'h7C;
                    16'h1A63: data_out = 8'h7D;
                    16'h1A64: data_out = 8'h7E;
                    16'h1A65: data_out = 8'h7F;
                    16'h1A66: data_out = 8'h80;
                    16'h1A67: data_out = 8'h81;
                    16'h1A68: data_out = 8'h82;
                    16'h1A69: data_out = 8'h83;
                    16'h1A6A: data_out = 8'h84;
                    16'h1A6B: data_out = 8'h85;
                    16'h1A6C: data_out = 8'h86;
                    16'h1A6D: data_out = 8'h87;
                    16'h1A6E: data_out = 8'h88;
                    16'h1A6F: data_out = 8'h89;
                    16'h1A70: data_out = 8'h8A;
                    16'h1A71: data_out = 8'h8B;
                    16'h1A72: data_out = 8'h8C;
                    16'h1A73: data_out = 8'h8D;
                    16'h1A74: data_out = 8'h8E;
                    16'h1A75: data_out = 8'h8F;
                    16'h1A76: data_out = 8'h90;
                    16'h1A77: data_out = 8'h91;
                    16'h1A78: data_out = 8'h92;
                    16'h1A79: data_out = 8'h93;
                    16'h1A7A: data_out = 8'h94;
                    16'h1A7B: data_out = 8'h95;
                    16'h1A7C: data_out = 8'h96;
                    16'h1A7D: data_out = 8'h97;
                    16'h1A7E: data_out = 8'h98;
                    16'h1A7F: data_out = 8'h99;
                    16'h1A80: data_out = 8'h1A;
                    16'h1A81: data_out = 8'h19;
                    16'h1A82: data_out = 8'h18;
                    16'h1A83: data_out = 8'h17;
                    16'h1A84: data_out = 8'h16;
                    16'h1A85: data_out = 8'h15;
                    16'h1A86: data_out = 8'h14;
                    16'h1A87: data_out = 8'h13;
                    16'h1A88: data_out = 8'h12;
                    16'h1A89: data_out = 8'h11;
                    16'h1A8A: data_out = 8'h10;
                    16'h1A8B: data_out = 8'hF;
                    16'h1A8C: data_out = 8'hE;
                    16'h1A8D: data_out = 8'hD;
                    16'h1A8E: data_out = 8'hC;
                    16'h1A8F: data_out = 8'hB;
                    16'h1A90: data_out = 8'hA;
                    16'h1A91: data_out = 8'h9;
                    16'h1A92: data_out = 8'h8;
                    16'h1A93: data_out = 8'h7;
                    16'h1A94: data_out = 8'h6;
                    16'h1A95: data_out = 8'h5;
                    16'h1A96: data_out = 8'h4;
                    16'h1A97: data_out = 8'h3;
                    16'h1A98: data_out = 8'h2;
                    16'h1A99: data_out = 8'h1;
                    16'h1A9A: data_out = 8'h0;
                    16'h1A9B: data_out = 8'h81;
                    16'h1A9C: data_out = 8'h82;
                    16'h1A9D: data_out = 8'h83;
                    16'h1A9E: data_out = 8'h84;
                    16'h1A9F: data_out = 8'h85;
                    16'h1AA0: data_out = 8'h86;
                    16'h1AA1: data_out = 8'h87;
                    16'h1AA2: data_out = 8'h88;
                    16'h1AA3: data_out = 8'h89;
                    16'h1AA4: data_out = 8'h8A;
                    16'h1AA5: data_out = 8'h8B;
                    16'h1AA6: data_out = 8'h8C;
                    16'h1AA7: data_out = 8'h8D;
                    16'h1AA8: data_out = 8'h8E;
                    16'h1AA9: data_out = 8'h8F;
                    16'h1AAA: data_out = 8'h90;
                    16'h1AAB: data_out = 8'h91;
                    16'h1AAC: data_out = 8'h92;
                    16'h1AAD: data_out = 8'h93;
                    16'h1AAE: data_out = 8'h94;
                    16'h1AAF: data_out = 8'h95;
                    16'h1AB0: data_out = 8'h96;
                    16'h1AB1: data_out = 8'h97;
                    16'h1AB2: data_out = 8'h98;
                    16'h1AB3: data_out = 8'h99;
                    16'h1AB4: data_out = 8'h9A;
                    16'h1AB5: data_out = 8'h9B;
                    16'h1AB6: data_out = 8'h9C;
                    16'h1AB7: data_out = 8'h9D;
                    16'h1AB8: data_out = 8'h9E;
                    16'h1AB9: data_out = 8'h9F;
                    16'h1ABA: data_out = 8'hA0;
                    16'h1ABB: data_out = 8'hA1;
                    16'h1ABC: data_out = 8'hA2;
                    16'h1ABD: data_out = 8'hA3;
                    16'h1ABE: data_out = 8'hA4;
                    16'h1ABF: data_out = 8'hA5;
                    16'h1AC0: data_out = 8'hA6;
                    16'h1AC1: data_out = 8'hA7;
                    16'h1AC2: data_out = 8'hA8;
                    16'h1AC3: data_out = 8'hA9;
                    16'h1AC4: data_out = 8'hAA;
                    16'h1AC5: data_out = 8'hAB;
                    16'h1AC6: data_out = 8'hAC;
                    16'h1AC7: data_out = 8'hAD;
                    16'h1AC8: data_out = 8'hAE;
                    16'h1AC9: data_out = 8'hAF;
                    16'h1ACA: data_out = 8'hB0;
                    16'h1ACB: data_out = 8'hB1;
                    16'h1ACC: data_out = 8'hB2;
                    16'h1ACD: data_out = 8'hB3;
                    16'h1ACE: data_out = 8'hB4;
                    16'h1ACF: data_out = 8'hB5;
                    16'h1AD0: data_out = 8'hB6;
                    16'h1AD1: data_out = 8'hB7;
                    16'h1AD2: data_out = 8'hB8;
                    16'h1AD3: data_out = 8'hB9;
                    16'h1AD4: data_out = 8'hBA;
                    16'h1AD5: data_out = 8'hBB;
                    16'h1AD6: data_out = 8'hBC;
                    16'h1AD7: data_out = 8'hBD;
                    16'h1AD8: data_out = 8'hBE;
                    16'h1AD9: data_out = 8'hBF;
                    16'h1ADA: data_out = 8'hC0;
                    16'h1ADB: data_out = 8'hC1;
                    16'h1ADC: data_out = 8'hC2;
                    16'h1ADD: data_out = 8'hC3;
                    16'h1ADE: data_out = 8'hC4;
                    16'h1ADF: data_out = 8'hC5;
                    16'h1AE0: data_out = 8'hC6;
                    16'h1AE1: data_out = 8'hC7;
                    16'h1AE2: data_out = 8'hC8;
                    16'h1AE3: data_out = 8'hC9;
                    16'h1AE4: data_out = 8'hCA;
                    16'h1AE5: data_out = 8'hCB;
                    16'h1AE6: data_out = 8'hCC;
                    16'h1AE7: data_out = 8'hCD;
                    16'h1AE8: data_out = 8'hCE;
                    16'h1AE9: data_out = 8'hCF;
                    16'h1AEA: data_out = 8'hD0;
                    16'h1AEB: data_out = 8'hD1;
                    16'h1AEC: data_out = 8'hD2;
                    16'h1AED: data_out = 8'hD3;
                    16'h1AEE: data_out = 8'hD4;
                    16'h1AEF: data_out = 8'hD5;
                    16'h1AF0: data_out = 8'hD6;
                    16'h1AF1: data_out = 8'hD7;
                    16'h1AF2: data_out = 8'hD8;
                    16'h1AF3: data_out = 8'hD9;
                    16'h1AF4: data_out = 8'hDA;
                    16'h1AF5: data_out = 8'hDB;
                    16'h1AF6: data_out = 8'hDC;
                    16'h1AF7: data_out = 8'hDD;
                    16'h1AF8: data_out = 8'hDE;
                    16'h1AF9: data_out = 8'hDF;
                    16'h1AFA: data_out = 8'hE0;
                    16'h1AFB: data_out = 8'hE1;
                    16'h1AFC: data_out = 8'hE2;
                    16'h1AFD: data_out = 8'hE3;
                    16'h1AFE: data_out = 8'hE4;
                    16'h1AFF: data_out = 8'hE5;
                    16'h1B00: data_out = 8'h1B;
                    16'h1B01: data_out = 8'h1C;
                    16'h1B02: data_out = 8'h1D;
                    16'h1B03: data_out = 8'h1E;
                    16'h1B04: data_out = 8'h1F;
                    16'h1B05: data_out = 8'h20;
                    16'h1B06: data_out = 8'h21;
                    16'h1B07: data_out = 8'h22;
                    16'h1B08: data_out = 8'h23;
                    16'h1B09: data_out = 8'h24;
                    16'h1B0A: data_out = 8'h25;
                    16'h1B0B: data_out = 8'h26;
                    16'h1B0C: data_out = 8'h27;
                    16'h1B0D: data_out = 8'h28;
                    16'h1B0E: data_out = 8'h29;
                    16'h1B0F: data_out = 8'h2A;
                    16'h1B10: data_out = 8'h2B;
                    16'h1B11: data_out = 8'h2C;
                    16'h1B12: data_out = 8'h2D;
                    16'h1B13: data_out = 8'h2E;
                    16'h1B14: data_out = 8'h2F;
                    16'h1B15: data_out = 8'h30;
                    16'h1B16: data_out = 8'h31;
                    16'h1B17: data_out = 8'h32;
                    16'h1B18: data_out = 8'h33;
                    16'h1B19: data_out = 8'h34;
                    16'h1B1A: data_out = 8'h35;
                    16'h1B1B: data_out = 8'h36;
                    16'h1B1C: data_out = 8'h37;
                    16'h1B1D: data_out = 8'h38;
                    16'h1B1E: data_out = 8'h39;
                    16'h1B1F: data_out = 8'h3A;
                    16'h1B20: data_out = 8'h3B;
                    16'h1B21: data_out = 8'h3C;
                    16'h1B22: data_out = 8'h3D;
                    16'h1B23: data_out = 8'h3E;
                    16'h1B24: data_out = 8'h3F;
                    16'h1B25: data_out = 8'h40;
                    16'h1B26: data_out = 8'h41;
                    16'h1B27: data_out = 8'h42;
                    16'h1B28: data_out = 8'h43;
                    16'h1B29: data_out = 8'h44;
                    16'h1B2A: data_out = 8'h45;
                    16'h1B2B: data_out = 8'h46;
                    16'h1B2C: data_out = 8'h47;
                    16'h1B2D: data_out = 8'h48;
                    16'h1B2E: data_out = 8'h49;
                    16'h1B2F: data_out = 8'h4A;
                    16'h1B30: data_out = 8'h4B;
                    16'h1B31: data_out = 8'h4C;
                    16'h1B32: data_out = 8'h4D;
                    16'h1B33: data_out = 8'h4E;
                    16'h1B34: data_out = 8'h4F;
                    16'h1B35: data_out = 8'h50;
                    16'h1B36: data_out = 8'h51;
                    16'h1B37: data_out = 8'h52;
                    16'h1B38: data_out = 8'h53;
                    16'h1B39: data_out = 8'h54;
                    16'h1B3A: data_out = 8'h55;
                    16'h1B3B: data_out = 8'h56;
                    16'h1B3C: data_out = 8'h57;
                    16'h1B3D: data_out = 8'h58;
                    16'h1B3E: data_out = 8'h59;
                    16'h1B3F: data_out = 8'h5A;
                    16'h1B40: data_out = 8'h5B;
                    16'h1B41: data_out = 8'h5C;
                    16'h1B42: data_out = 8'h5D;
                    16'h1B43: data_out = 8'h5E;
                    16'h1B44: data_out = 8'h5F;
                    16'h1B45: data_out = 8'h60;
                    16'h1B46: data_out = 8'h61;
                    16'h1B47: data_out = 8'h62;
                    16'h1B48: data_out = 8'h63;
                    16'h1B49: data_out = 8'h64;
                    16'h1B4A: data_out = 8'h65;
                    16'h1B4B: data_out = 8'h66;
                    16'h1B4C: data_out = 8'h67;
                    16'h1B4D: data_out = 8'h68;
                    16'h1B4E: data_out = 8'h69;
                    16'h1B4F: data_out = 8'h6A;
                    16'h1B50: data_out = 8'h6B;
                    16'h1B51: data_out = 8'h6C;
                    16'h1B52: data_out = 8'h6D;
                    16'h1B53: data_out = 8'h6E;
                    16'h1B54: data_out = 8'h6F;
                    16'h1B55: data_out = 8'h70;
                    16'h1B56: data_out = 8'h71;
                    16'h1B57: data_out = 8'h72;
                    16'h1B58: data_out = 8'h73;
                    16'h1B59: data_out = 8'h74;
                    16'h1B5A: data_out = 8'h75;
                    16'h1B5B: data_out = 8'h76;
                    16'h1B5C: data_out = 8'h77;
                    16'h1B5D: data_out = 8'h78;
                    16'h1B5E: data_out = 8'h79;
                    16'h1B5F: data_out = 8'h7A;
                    16'h1B60: data_out = 8'h7B;
                    16'h1B61: data_out = 8'h7C;
                    16'h1B62: data_out = 8'h7D;
                    16'h1B63: data_out = 8'h7E;
                    16'h1B64: data_out = 8'h7F;
                    16'h1B65: data_out = 8'h80;
                    16'h1B66: data_out = 8'h81;
                    16'h1B67: data_out = 8'h82;
                    16'h1B68: data_out = 8'h83;
                    16'h1B69: data_out = 8'h84;
                    16'h1B6A: data_out = 8'h85;
                    16'h1B6B: data_out = 8'h86;
                    16'h1B6C: data_out = 8'h87;
                    16'h1B6D: data_out = 8'h88;
                    16'h1B6E: data_out = 8'h89;
                    16'h1B6F: data_out = 8'h8A;
                    16'h1B70: data_out = 8'h8B;
                    16'h1B71: data_out = 8'h8C;
                    16'h1B72: data_out = 8'h8D;
                    16'h1B73: data_out = 8'h8E;
                    16'h1B74: data_out = 8'h8F;
                    16'h1B75: data_out = 8'h90;
                    16'h1B76: data_out = 8'h91;
                    16'h1B77: data_out = 8'h92;
                    16'h1B78: data_out = 8'h93;
                    16'h1B79: data_out = 8'h94;
                    16'h1B7A: data_out = 8'h95;
                    16'h1B7B: data_out = 8'h96;
                    16'h1B7C: data_out = 8'h97;
                    16'h1B7D: data_out = 8'h98;
                    16'h1B7E: data_out = 8'h99;
                    16'h1B7F: data_out = 8'h9A;
                    16'h1B80: data_out = 8'h1B;
                    16'h1B81: data_out = 8'h1A;
                    16'h1B82: data_out = 8'h19;
                    16'h1B83: data_out = 8'h18;
                    16'h1B84: data_out = 8'h17;
                    16'h1B85: data_out = 8'h16;
                    16'h1B86: data_out = 8'h15;
                    16'h1B87: data_out = 8'h14;
                    16'h1B88: data_out = 8'h13;
                    16'h1B89: data_out = 8'h12;
                    16'h1B8A: data_out = 8'h11;
                    16'h1B8B: data_out = 8'h10;
                    16'h1B8C: data_out = 8'hF;
                    16'h1B8D: data_out = 8'hE;
                    16'h1B8E: data_out = 8'hD;
                    16'h1B8F: data_out = 8'hC;
                    16'h1B90: data_out = 8'hB;
                    16'h1B91: data_out = 8'hA;
                    16'h1B92: data_out = 8'h9;
                    16'h1B93: data_out = 8'h8;
                    16'h1B94: data_out = 8'h7;
                    16'h1B95: data_out = 8'h6;
                    16'h1B96: data_out = 8'h5;
                    16'h1B97: data_out = 8'h4;
                    16'h1B98: data_out = 8'h3;
                    16'h1B99: data_out = 8'h2;
                    16'h1B9A: data_out = 8'h1;
                    16'h1B9B: data_out = 8'h0;
                    16'h1B9C: data_out = 8'h81;
                    16'h1B9D: data_out = 8'h82;
                    16'h1B9E: data_out = 8'h83;
                    16'h1B9F: data_out = 8'h84;
                    16'h1BA0: data_out = 8'h85;
                    16'h1BA1: data_out = 8'h86;
                    16'h1BA2: data_out = 8'h87;
                    16'h1BA3: data_out = 8'h88;
                    16'h1BA4: data_out = 8'h89;
                    16'h1BA5: data_out = 8'h8A;
                    16'h1BA6: data_out = 8'h8B;
                    16'h1BA7: data_out = 8'h8C;
                    16'h1BA8: data_out = 8'h8D;
                    16'h1BA9: data_out = 8'h8E;
                    16'h1BAA: data_out = 8'h8F;
                    16'h1BAB: data_out = 8'h90;
                    16'h1BAC: data_out = 8'h91;
                    16'h1BAD: data_out = 8'h92;
                    16'h1BAE: data_out = 8'h93;
                    16'h1BAF: data_out = 8'h94;
                    16'h1BB0: data_out = 8'h95;
                    16'h1BB1: data_out = 8'h96;
                    16'h1BB2: data_out = 8'h97;
                    16'h1BB3: data_out = 8'h98;
                    16'h1BB4: data_out = 8'h99;
                    16'h1BB5: data_out = 8'h9A;
                    16'h1BB6: data_out = 8'h9B;
                    16'h1BB7: data_out = 8'h9C;
                    16'h1BB8: data_out = 8'h9D;
                    16'h1BB9: data_out = 8'h9E;
                    16'h1BBA: data_out = 8'h9F;
                    16'h1BBB: data_out = 8'hA0;
                    16'h1BBC: data_out = 8'hA1;
                    16'h1BBD: data_out = 8'hA2;
                    16'h1BBE: data_out = 8'hA3;
                    16'h1BBF: data_out = 8'hA4;
                    16'h1BC0: data_out = 8'hA5;
                    16'h1BC1: data_out = 8'hA6;
                    16'h1BC2: data_out = 8'hA7;
                    16'h1BC3: data_out = 8'hA8;
                    16'h1BC4: data_out = 8'hA9;
                    16'h1BC5: data_out = 8'hAA;
                    16'h1BC6: data_out = 8'hAB;
                    16'h1BC7: data_out = 8'hAC;
                    16'h1BC8: data_out = 8'hAD;
                    16'h1BC9: data_out = 8'hAE;
                    16'h1BCA: data_out = 8'hAF;
                    16'h1BCB: data_out = 8'hB0;
                    16'h1BCC: data_out = 8'hB1;
                    16'h1BCD: data_out = 8'hB2;
                    16'h1BCE: data_out = 8'hB3;
                    16'h1BCF: data_out = 8'hB4;
                    16'h1BD0: data_out = 8'hB5;
                    16'h1BD1: data_out = 8'hB6;
                    16'h1BD2: data_out = 8'hB7;
                    16'h1BD3: data_out = 8'hB8;
                    16'h1BD4: data_out = 8'hB9;
                    16'h1BD5: data_out = 8'hBA;
                    16'h1BD6: data_out = 8'hBB;
                    16'h1BD7: data_out = 8'hBC;
                    16'h1BD8: data_out = 8'hBD;
                    16'h1BD9: data_out = 8'hBE;
                    16'h1BDA: data_out = 8'hBF;
                    16'h1BDB: data_out = 8'hC0;
                    16'h1BDC: data_out = 8'hC1;
                    16'h1BDD: data_out = 8'hC2;
                    16'h1BDE: data_out = 8'hC3;
                    16'h1BDF: data_out = 8'hC4;
                    16'h1BE0: data_out = 8'hC5;
                    16'h1BE1: data_out = 8'hC6;
                    16'h1BE2: data_out = 8'hC7;
                    16'h1BE3: data_out = 8'hC8;
                    16'h1BE4: data_out = 8'hC9;
                    16'h1BE5: data_out = 8'hCA;
                    16'h1BE6: data_out = 8'hCB;
                    16'h1BE7: data_out = 8'hCC;
                    16'h1BE8: data_out = 8'hCD;
                    16'h1BE9: data_out = 8'hCE;
                    16'h1BEA: data_out = 8'hCF;
                    16'h1BEB: data_out = 8'hD0;
                    16'h1BEC: data_out = 8'hD1;
                    16'h1BED: data_out = 8'hD2;
                    16'h1BEE: data_out = 8'hD3;
                    16'h1BEF: data_out = 8'hD4;
                    16'h1BF0: data_out = 8'hD5;
                    16'h1BF1: data_out = 8'hD6;
                    16'h1BF2: data_out = 8'hD7;
                    16'h1BF3: data_out = 8'hD8;
                    16'h1BF4: data_out = 8'hD9;
                    16'h1BF5: data_out = 8'hDA;
                    16'h1BF6: data_out = 8'hDB;
                    16'h1BF7: data_out = 8'hDC;
                    16'h1BF8: data_out = 8'hDD;
                    16'h1BF9: data_out = 8'hDE;
                    16'h1BFA: data_out = 8'hDF;
                    16'h1BFB: data_out = 8'hE0;
                    16'h1BFC: data_out = 8'hE1;
                    16'h1BFD: data_out = 8'hE2;
                    16'h1BFE: data_out = 8'hE3;
                    16'h1BFF: data_out = 8'hE4;
                    16'h1C00: data_out = 8'h1C;
                    16'h1C01: data_out = 8'h1D;
                    16'h1C02: data_out = 8'h1E;
                    16'h1C03: data_out = 8'h1F;
                    16'h1C04: data_out = 8'h20;
                    16'h1C05: data_out = 8'h21;
                    16'h1C06: data_out = 8'h22;
                    16'h1C07: data_out = 8'h23;
                    16'h1C08: data_out = 8'h24;
                    16'h1C09: data_out = 8'h25;
                    16'h1C0A: data_out = 8'h26;
                    16'h1C0B: data_out = 8'h27;
                    16'h1C0C: data_out = 8'h28;
                    16'h1C0D: data_out = 8'h29;
                    16'h1C0E: data_out = 8'h2A;
                    16'h1C0F: data_out = 8'h2B;
                    16'h1C10: data_out = 8'h2C;
                    16'h1C11: data_out = 8'h2D;
                    16'h1C12: data_out = 8'h2E;
                    16'h1C13: data_out = 8'h2F;
                    16'h1C14: data_out = 8'h30;
                    16'h1C15: data_out = 8'h31;
                    16'h1C16: data_out = 8'h32;
                    16'h1C17: data_out = 8'h33;
                    16'h1C18: data_out = 8'h34;
                    16'h1C19: data_out = 8'h35;
                    16'h1C1A: data_out = 8'h36;
                    16'h1C1B: data_out = 8'h37;
                    16'h1C1C: data_out = 8'h38;
                    16'h1C1D: data_out = 8'h39;
                    16'h1C1E: data_out = 8'h3A;
                    16'h1C1F: data_out = 8'h3B;
                    16'h1C20: data_out = 8'h3C;
                    16'h1C21: data_out = 8'h3D;
                    16'h1C22: data_out = 8'h3E;
                    16'h1C23: data_out = 8'h3F;
                    16'h1C24: data_out = 8'h40;
                    16'h1C25: data_out = 8'h41;
                    16'h1C26: data_out = 8'h42;
                    16'h1C27: data_out = 8'h43;
                    16'h1C28: data_out = 8'h44;
                    16'h1C29: data_out = 8'h45;
                    16'h1C2A: data_out = 8'h46;
                    16'h1C2B: data_out = 8'h47;
                    16'h1C2C: data_out = 8'h48;
                    16'h1C2D: data_out = 8'h49;
                    16'h1C2E: data_out = 8'h4A;
                    16'h1C2F: data_out = 8'h4B;
                    16'h1C30: data_out = 8'h4C;
                    16'h1C31: data_out = 8'h4D;
                    16'h1C32: data_out = 8'h4E;
                    16'h1C33: data_out = 8'h4F;
                    16'h1C34: data_out = 8'h50;
                    16'h1C35: data_out = 8'h51;
                    16'h1C36: data_out = 8'h52;
                    16'h1C37: data_out = 8'h53;
                    16'h1C38: data_out = 8'h54;
                    16'h1C39: data_out = 8'h55;
                    16'h1C3A: data_out = 8'h56;
                    16'h1C3B: data_out = 8'h57;
                    16'h1C3C: data_out = 8'h58;
                    16'h1C3D: data_out = 8'h59;
                    16'h1C3E: data_out = 8'h5A;
                    16'h1C3F: data_out = 8'h5B;
                    16'h1C40: data_out = 8'h5C;
                    16'h1C41: data_out = 8'h5D;
                    16'h1C42: data_out = 8'h5E;
                    16'h1C43: data_out = 8'h5F;
                    16'h1C44: data_out = 8'h60;
                    16'h1C45: data_out = 8'h61;
                    16'h1C46: data_out = 8'h62;
                    16'h1C47: data_out = 8'h63;
                    16'h1C48: data_out = 8'h64;
                    16'h1C49: data_out = 8'h65;
                    16'h1C4A: data_out = 8'h66;
                    16'h1C4B: data_out = 8'h67;
                    16'h1C4C: data_out = 8'h68;
                    16'h1C4D: data_out = 8'h69;
                    16'h1C4E: data_out = 8'h6A;
                    16'h1C4F: data_out = 8'h6B;
                    16'h1C50: data_out = 8'h6C;
                    16'h1C51: data_out = 8'h6D;
                    16'h1C52: data_out = 8'h6E;
                    16'h1C53: data_out = 8'h6F;
                    16'h1C54: data_out = 8'h70;
                    16'h1C55: data_out = 8'h71;
                    16'h1C56: data_out = 8'h72;
                    16'h1C57: data_out = 8'h73;
                    16'h1C58: data_out = 8'h74;
                    16'h1C59: data_out = 8'h75;
                    16'h1C5A: data_out = 8'h76;
                    16'h1C5B: data_out = 8'h77;
                    16'h1C5C: data_out = 8'h78;
                    16'h1C5D: data_out = 8'h79;
                    16'h1C5E: data_out = 8'h7A;
                    16'h1C5F: data_out = 8'h7B;
                    16'h1C60: data_out = 8'h7C;
                    16'h1C61: data_out = 8'h7D;
                    16'h1C62: data_out = 8'h7E;
                    16'h1C63: data_out = 8'h7F;
                    16'h1C64: data_out = 8'h80;
                    16'h1C65: data_out = 8'h81;
                    16'h1C66: data_out = 8'h82;
                    16'h1C67: data_out = 8'h83;
                    16'h1C68: data_out = 8'h84;
                    16'h1C69: data_out = 8'h85;
                    16'h1C6A: data_out = 8'h86;
                    16'h1C6B: data_out = 8'h87;
                    16'h1C6C: data_out = 8'h88;
                    16'h1C6D: data_out = 8'h89;
                    16'h1C6E: data_out = 8'h8A;
                    16'h1C6F: data_out = 8'h8B;
                    16'h1C70: data_out = 8'h8C;
                    16'h1C71: data_out = 8'h8D;
                    16'h1C72: data_out = 8'h8E;
                    16'h1C73: data_out = 8'h8F;
                    16'h1C74: data_out = 8'h90;
                    16'h1C75: data_out = 8'h91;
                    16'h1C76: data_out = 8'h92;
                    16'h1C77: data_out = 8'h93;
                    16'h1C78: data_out = 8'h94;
                    16'h1C79: data_out = 8'h95;
                    16'h1C7A: data_out = 8'h96;
                    16'h1C7B: data_out = 8'h97;
                    16'h1C7C: data_out = 8'h98;
                    16'h1C7D: data_out = 8'h99;
                    16'h1C7E: data_out = 8'h9A;
                    16'h1C7F: data_out = 8'h9B;
                    16'h1C80: data_out = 8'h1C;
                    16'h1C81: data_out = 8'h1B;
                    16'h1C82: data_out = 8'h1A;
                    16'h1C83: data_out = 8'h19;
                    16'h1C84: data_out = 8'h18;
                    16'h1C85: data_out = 8'h17;
                    16'h1C86: data_out = 8'h16;
                    16'h1C87: data_out = 8'h15;
                    16'h1C88: data_out = 8'h14;
                    16'h1C89: data_out = 8'h13;
                    16'h1C8A: data_out = 8'h12;
                    16'h1C8B: data_out = 8'h11;
                    16'h1C8C: data_out = 8'h10;
                    16'h1C8D: data_out = 8'hF;
                    16'h1C8E: data_out = 8'hE;
                    16'h1C8F: data_out = 8'hD;
                    16'h1C90: data_out = 8'hC;
                    16'h1C91: data_out = 8'hB;
                    16'h1C92: data_out = 8'hA;
                    16'h1C93: data_out = 8'h9;
                    16'h1C94: data_out = 8'h8;
                    16'h1C95: data_out = 8'h7;
                    16'h1C96: data_out = 8'h6;
                    16'h1C97: data_out = 8'h5;
                    16'h1C98: data_out = 8'h4;
                    16'h1C99: data_out = 8'h3;
                    16'h1C9A: data_out = 8'h2;
                    16'h1C9B: data_out = 8'h1;
                    16'h1C9C: data_out = 8'h0;
                    16'h1C9D: data_out = 8'h81;
                    16'h1C9E: data_out = 8'h82;
                    16'h1C9F: data_out = 8'h83;
                    16'h1CA0: data_out = 8'h84;
                    16'h1CA1: data_out = 8'h85;
                    16'h1CA2: data_out = 8'h86;
                    16'h1CA3: data_out = 8'h87;
                    16'h1CA4: data_out = 8'h88;
                    16'h1CA5: data_out = 8'h89;
                    16'h1CA6: data_out = 8'h8A;
                    16'h1CA7: data_out = 8'h8B;
                    16'h1CA8: data_out = 8'h8C;
                    16'h1CA9: data_out = 8'h8D;
                    16'h1CAA: data_out = 8'h8E;
                    16'h1CAB: data_out = 8'h8F;
                    16'h1CAC: data_out = 8'h90;
                    16'h1CAD: data_out = 8'h91;
                    16'h1CAE: data_out = 8'h92;
                    16'h1CAF: data_out = 8'h93;
                    16'h1CB0: data_out = 8'h94;
                    16'h1CB1: data_out = 8'h95;
                    16'h1CB2: data_out = 8'h96;
                    16'h1CB3: data_out = 8'h97;
                    16'h1CB4: data_out = 8'h98;
                    16'h1CB5: data_out = 8'h99;
                    16'h1CB6: data_out = 8'h9A;
                    16'h1CB7: data_out = 8'h9B;
                    16'h1CB8: data_out = 8'h9C;
                    16'h1CB9: data_out = 8'h9D;
                    16'h1CBA: data_out = 8'h9E;
                    16'h1CBB: data_out = 8'h9F;
                    16'h1CBC: data_out = 8'hA0;
                    16'h1CBD: data_out = 8'hA1;
                    16'h1CBE: data_out = 8'hA2;
                    16'h1CBF: data_out = 8'hA3;
                    16'h1CC0: data_out = 8'hA4;
                    16'h1CC1: data_out = 8'hA5;
                    16'h1CC2: data_out = 8'hA6;
                    16'h1CC3: data_out = 8'hA7;
                    16'h1CC4: data_out = 8'hA8;
                    16'h1CC5: data_out = 8'hA9;
                    16'h1CC6: data_out = 8'hAA;
                    16'h1CC7: data_out = 8'hAB;
                    16'h1CC8: data_out = 8'hAC;
                    16'h1CC9: data_out = 8'hAD;
                    16'h1CCA: data_out = 8'hAE;
                    16'h1CCB: data_out = 8'hAF;
                    16'h1CCC: data_out = 8'hB0;
                    16'h1CCD: data_out = 8'hB1;
                    16'h1CCE: data_out = 8'hB2;
                    16'h1CCF: data_out = 8'hB3;
                    16'h1CD0: data_out = 8'hB4;
                    16'h1CD1: data_out = 8'hB5;
                    16'h1CD2: data_out = 8'hB6;
                    16'h1CD3: data_out = 8'hB7;
                    16'h1CD4: data_out = 8'hB8;
                    16'h1CD5: data_out = 8'hB9;
                    16'h1CD6: data_out = 8'hBA;
                    16'h1CD7: data_out = 8'hBB;
                    16'h1CD8: data_out = 8'hBC;
                    16'h1CD9: data_out = 8'hBD;
                    16'h1CDA: data_out = 8'hBE;
                    16'h1CDB: data_out = 8'hBF;
                    16'h1CDC: data_out = 8'hC0;
                    16'h1CDD: data_out = 8'hC1;
                    16'h1CDE: data_out = 8'hC2;
                    16'h1CDF: data_out = 8'hC3;
                    16'h1CE0: data_out = 8'hC4;
                    16'h1CE1: data_out = 8'hC5;
                    16'h1CE2: data_out = 8'hC6;
                    16'h1CE3: data_out = 8'hC7;
                    16'h1CE4: data_out = 8'hC8;
                    16'h1CE5: data_out = 8'hC9;
                    16'h1CE6: data_out = 8'hCA;
                    16'h1CE7: data_out = 8'hCB;
                    16'h1CE8: data_out = 8'hCC;
                    16'h1CE9: data_out = 8'hCD;
                    16'h1CEA: data_out = 8'hCE;
                    16'h1CEB: data_out = 8'hCF;
                    16'h1CEC: data_out = 8'hD0;
                    16'h1CED: data_out = 8'hD1;
                    16'h1CEE: data_out = 8'hD2;
                    16'h1CEF: data_out = 8'hD3;
                    16'h1CF0: data_out = 8'hD4;
                    16'h1CF1: data_out = 8'hD5;
                    16'h1CF2: data_out = 8'hD6;
                    16'h1CF3: data_out = 8'hD7;
                    16'h1CF4: data_out = 8'hD8;
                    16'h1CF5: data_out = 8'hD9;
                    16'h1CF6: data_out = 8'hDA;
                    16'h1CF7: data_out = 8'hDB;
                    16'h1CF8: data_out = 8'hDC;
                    16'h1CF9: data_out = 8'hDD;
                    16'h1CFA: data_out = 8'hDE;
                    16'h1CFB: data_out = 8'hDF;
                    16'h1CFC: data_out = 8'hE0;
                    16'h1CFD: data_out = 8'hE1;
                    16'h1CFE: data_out = 8'hE2;
                    16'h1CFF: data_out = 8'hE3;
                    16'h1D00: data_out = 8'h1D;
                    16'h1D01: data_out = 8'h1E;
                    16'h1D02: data_out = 8'h1F;
                    16'h1D03: data_out = 8'h20;
                    16'h1D04: data_out = 8'h21;
                    16'h1D05: data_out = 8'h22;
                    16'h1D06: data_out = 8'h23;
                    16'h1D07: data_out = 8'h24;
                    16'h1D08: data_out = 8'h25;
                    16'h1D09: data_out = 8'h26;
                    16'h1D0A: data_out = 8'h27;
                    16'h1D0B: data_out = 8'h28;
                    16'h1D0C: data_out = 8'h29;
                    16'h1D0D: data_out = 8'h2A;
                    16'h1D0E: data_out = 8'h2B;
                    16'h1D0F: data_out = 8'h2C;
                    16'h1D10: data_out = 8'h2D;
                    16'h1D11: data_out = 8'h2E;
                    16'h1D12: data_out = 8'h2F;
                    16'h1D13: data_out = 8'h30;
                    16'h1D14: data_out = 8'h31;
                    16'h1D15: data_out = 8'h32;
                    16'h1D16: data_out = 8'h33;
                    16'h1D17: data_out = 8'h34;
                    16'h1D18: data_out = 8'h35;
                    16'h1D19: data_out = 8'h36;
                    16'h1D1A: data_out = 8'h37;
                    16'h1D1B: data_out = 8'h38;
                    16'h1D1C: data_out = 8'h39;
                    16'h1D1D: data_out = 8'h3A;
                    16'h1D1E: data_out = 8'h3B;
                    16'h1D1F: data_out = 8'h3C;
                    16'h1D20: data_out = 8'h3D;
                    16'h1D21: data_out = 8'h3E;
                    16'h1D22: data_out = 8'h3F;
                    16'h1D23: data_out = 8'h40;
                    16'h1D24: data_out = 8'h41;
                    16'h1D25: data_out = 8'h42;
                    16'h1D26: data_out = 8'h43;
                    16'h1D27: data_out = 8'h44;
                    16'h1D28: data_out = 8'h45;
                    16'h1D29: data_out = 8'h46;
                    16'h1D2A: data_out = 8'h47;
                    16'h1D2B: data_out = 8'h48;
                    16'h1D2C: data_out = 8'h49;
                    16'h1D2D: data_out = 8'h4A;
                    16'h1D2E: data_out = 8'h4B;
                    16'h1D2F: data_out = 8'h4C;
                    16'h1D30: data_out = 8'h4D;
                    16'h1D31: data_out = 8'h4E;
                    16'h1D32: data_out = 8'h4F;
                    16'h1D33: data_out = 8'h50;
                    16'h1D34: data_out = 8'h51;
                    16'h1D35: data_out = 8'h52;
                    16'h1D36: data_out = 8'h53;
                    16'h1D37: data_out = 8'h54;
                    16'h1D38: data_out = 8'h55;
                    16'h1D39: data_out = 8'h56;
                    16'h1D3A: data_out = 8'h57;
                    16'h1D3B: data_out = 8'h58;
                    16'h1D3C: data_out = 8'h59;
                    16'h1D3D: data_out = 8'h5A;
                    16'h1D3E: data_out = 8'h5B;
                    16'h1D3F: data_out = 8'h5C;
                    16'h1D40: data_out = 8'h5D;
                    16'h1D41: data_out = 8'h5E;
                    16'h1D42: data_out = 8'h5F;
                    16'h1D43: data_out = 8'h60;
                    16'h1D44: data_out = 8'h61;
                    16'h1D45: data_out = 8'h62;
                    16'h1D46: data_out = 8'h63;
                    16'h1D47: data_out = 8'h64;
                    16'h1D48: data_out = 8'h65;
                    16'h1D49: data_out = 8'h66;
                    16'h1D4A: data_out = 8'h67;
                    16'h1D4B: data_out = 8'h68;
                    16'h1D4C: data_out = 8'h69;
                    16'h1D4D: data_out = 8'h6A;
                    16'h1D4E: data_out = 8'h6B;
                    16'h1D4F: data_out = 8'h6C;
                    16'h1D50: data_out = 8'h6D;
                    16'h1D51: data_out = 8'h6E;
                    16'h1D52: data_out = 8'h6F;
                    16'h1D53: data_out = 8'h70;
                    16'h1D54: data_out = 8'h71;
                    16'h1D55: data_out = 8'h72;
                    16'h1D56: data_out = 8'h73;
                    16'h1D57: data_out = 8'h74;
                    16'h1D58: data_out = 8'h75;
                    16'h1D59: data_out = 8'h76;
                    16'h1D5A: data_out = 8'h77;
                    16'h1D5B: data_out = 8'h78;
                    16'h1D5C: data_out = 8'h79;
                    16'h1D5D: data_out = 8'h7A;
                    16'h1D5E: data_out = 8'h7B;
                    16'h1D5F: data_out = 8'h7C;
                    16'h1D60: data_out = 8'h7D;
                    16'h1D61: data_out = 8'h7E;
                    16'h1D62: data_out = 8'h7F;
                    16'h1D63: data_out = 8'h80;
                    16'h1D64: data_out = 8'h81;
                    16'h1D65: data_out = 8'h82;
                    16'h1D66: data_out = 8'h83;
                    16'h1D67: data_out = 8'h84;
                    16'h1D68: data_out = 8'h85;
                    16'h1D69: data_out = 8'h86;
                    16'h1D6A: data_out = 8'h87;
                    16'h1D6B: data_out = 8'h88;
                    16'h1D6C: data_out = 8'h89;
                    16'h1D6D: data_out = 8'h8A;
                    16'h1D6E: data_out = 8'h8B;
                    16'h1D6F: data_out = 8'h8C;
                    16'h1D70: data_out = 8'h8D;
                    16'h1D71: data_out = 8'h8E;
                    16'h1D72: data_out = 8'h8F;
                    16'h1D73: data_out = 8'h90;
                    16'h1D74: data_out = 8'h91;
                    16'h1D75: data_out = 8'h92;
                    16'h1D76: data_out = 8'h93;
                    16'h1D77: data_out = 8'h94;
                    16'h1D78: data_out = 8'h95;
                    16'h1D79: data_out = 8'h96;
                    16'h1D7A: data_out = 8'h97;
                    16'h1D7B: data_out = 8'h98;
                    16'h1D7C: data_out = 8'h99;
                    16'h1D7D: data_out = 8'h9A;
                    16'h1D7E: data_out = 8'h9B;
                    16'h1D7F: data_out = 8'h9C;
                    16'h1D80: data_out = 8'h1D;
                    16'h1D81: data_out = 8'h1C;
                    16'h1D82: data_out = 8'h1B;
                    16'h1D83: data_out = 8'h1A;
                    16'h1D84: data_out = 8'h19;
                    16'h1D85: data_out = 8'h18;
                    16'h1D86: data_out = 8'h17;
                    16'h1D87: data_out = 8'h16;
                    16'h1D88: data_out = 8'h15;
                    16'h1D89: data_out = 8'h14;
                    16'h1D8A: data_out = 8'h13;
                    16'h1D8B: data_out = 8'h12;
                    16'h1D8C: data_out = 8'h11;
                    16'h1D8D: data_out = 8'h10;
                    16'h1D8E: data_out = 8'hF;
                    16'h1D8F: data_out = 8'hE;
                    16'h1D90: data_out = 8'hD;
                    16'h1D91: data_out = 8'hC;
                    16'h1D92: data_out = 8'hB;
                    16'h1D93: data_out = 8'hA;
                    16'h1D94: data_out = 8'h9;
                    16'h1D95: data_out = 8'h8;
                    16'h1D96: data_out = 8'h7;
                    16'h1D97: data_out = 8'h6;
                    16'h1D98: data_out = 8'h5;
                    16'h1D99: data_out = 8'h4;
                    16'h1D9A: data_out = 8'h3;
                    16'h1D9B: data_out = 8'h2;
                    16'h1D9C: data_out = 8'h1;
                    16'h1D9D: data_out = 8'h0;
                    16'h1D9E: data_out = 8'h81;
                    16'h1D9F: data_out = 8'h82;
                    16'h1DA0: data_out = 8'h83;
                    16'h1DA1: data_out = 8'h84;
                    16'h1DA2: data_out = 8'h85;
                    16'h1DA3: data_out = 8'h86;
                    16'h1DA4: data_out = 8'h87;
                    16'h1DA5: data_out = 8'h88;
                    16'h1DA6: data_out = 8'h89;
                    16'h1DA7: data_out = 8'h8A;
                    16'h1DA8: data_out = 8'h8B;
                    16'h1DA9: data_out = 8'h8C;
                    16'h1DAA: data_out = 8'h8D;
                    16'h1DAB: data_out = 8'h8E;
                    16'h1DAC: data_out = 8'h8F;
                    16'h1DAD: data_out = 8'h90;
                    16'h1DAE: data_out = 8'h91;
                    16'h1DAF: data_out = 8'h92;
                    16'h1DB0: data_out = 8'h93;
                    16'h1DB1: data_out = 8'h94;
                    16'h1DB2: data_out = 8'h95;
                    16'h1DB3: data_out = 8'h96;
                    16'h1DB4: data_out = 8'h97;
                    16'h1DB5: data_out = 8'h98;
                    16'h1DB6: data_out = 8'h99;
                    16'h1DB7: data_out = 8'h9A;
                    16'h1DB8: data_out = 8'h9B;
                    16'h1DB9: data_out = 8'h9C;
                    16'h1DBA: data_out = 8'h9D;
                    16'h1DBB: data_out = 8'h9E;
                    16'h1DBC: data_out = 8'h9F;
                    16'h1DBD: data_out = 8'hA0;
                    16'h1DBE: data_out = 8'hA1;
                    16'h1DBF: data_out = 8'hA2;
                    16'h1DC0: data_out = 8'hA3;
                    16'h1DC1: data_out = 8'hA4;
                    16'h1DC2: data_out = 8'hA5;
                    16'h1DC3: data_out = 8'hA6;
                    16'h1DC4: data_out = 8'hA7;
                    16'h1DC5: data_out = 8'hA8;
                    16'h1DC6: data_out = 8'hA9;
                    16'h1DC7: data_out = 8'hAA;
                    16'h1DC8: data_out = 8'hAB;
                    16'h1DC9: data_out = 8'hAC;
                    16'h1DCA: data_out = 8'hAD;
                    16'h1DCB: data_out = 8'hAE;
                    16'h1DCC: data_out = 8'hAF;
                    16'h1DCD: data_out = 8'hB0;
                    16'h1DCE: data_out = 8'hB1;
                    16'h1DCF: data_out = 8'hB2;
                    16'h1DD0: data_out = 8'hB3;
                    16'h1DD1: data_out = 8'hB4;
                    16'h1DD2: data_out = 8'hB5;
                    16'h1DD3: data_out = 8'hB6;
                    16'h1DD4: data_out = 8'hB7;
                    16'h1DD5: data_out = 8'hB8;
                    16'h1DD6: data_out = 8'hB9;
                    16'h1DD7: data_out = 8'hBA;
                    16'h1DD8: data_out = 8'hBB;
                    16'h1DD9: data_out = 8'hBC;
                    16'h1DDA: data_out = 8'hBD;
                    16'h1DDB: data_out = 8'hBE;
                    16'h1DDC: data_out = 8'hBF;
                    16'h1DDD: data_out = 8'hC0;
                    16'h1DDE: data_out = 8'hC1;
                    16'h1DDF: data_out = 8'hC2;
                    16'h1DE0: data_out = 8'hC3;
                    16'h1DE1: data_out = 8'hC4;
                    16'h1DE2: data_out = 8'hC5;
                    16'h1DE3: data_out = 8'hC6;
                    16'h1DE4: data_out = 8'hC7;
                    16'h1DE5: data_out = 8'hC8;
                    16'h1DE6: data_out = 8'hC9;
                    16'h1DE7: data_out = 8'hCA;
                    16'h1DE8: data_out = 8'hCB;
                    16'h1DE9: data_out = 8'hCC;
                    16'h1DEA: data_out = 8'hCD;
                    16'h1DEB: data_out = 8'hCE;
                    16'h1DEC: data_out = 8'hCF;
                    16'h1DED: data_out = 8'hD0;
                    16'h1DEE: data_out = 8'hD1;
                    16'h1DEF: data_out = 8'hD2;
                    16'h1DF0: data_out = 8'hD3;
                    16'h1DF1: data_out = 8'hD4;
                    16'h1DF2: data_out = 8'hD5;
                    16'h1DF3: data_out = 8'hD6;
                    16'h1DF4: data_out = 8'hD7;
                    16'h1DF5: data_out = 8'hD8;
                    16'h1DF6: data_out = 8'hD9;
                    16'h1DF7: data_out = 8'hDA;
                    16'h1DF8: data_out = 8'hDB;
                    16'h1DF9: data_out = 8'hDC;
                    16'h1DFA: data_out = 8'hDD;
                    16'h1DFB: data_out = 8'hDE;
                    16'h1DFC: data_out = 8'hDF;
                    16'h1DFD: data_out = 8'hE0;
                    16'h1DFE: data_out = 8'hE1;
                    16'h1DFF: data_out = 8'hE2;
                    16'h1E00: data_out = 8'h1E;
                    16'h1E01: data_out = 8'h1F;
                    16'h1E02: data_out = 8'h20;
                    16'h1E03: data_out = 8'h21;
                    16'h1E04: data_out = 8'h22;
                    16'h1E05: data_out = 8'h23;
                    16'h1E06: data_out = 8'h24;
                    16'h1E07: data_out = 8'h25;
                    16'h1E08: data_out = 8'h26;
                    16'h1E09: data_out = 8'h27;
                    16'h1E0A: data_out = 8'h28;
                    16'h1E0B: data_out = 8'h29;
                    16'h1E0C: data_out = 8'h2A;
                    16'h1E0D: data_out = 8'h2B;
                    16'h1E0E: data_out = 8'h2C;
                    16'h1E0F: data_out = 8'h2D;
                    16'h1E10: data_out = 8'h2E;
                    16'h1E11: data_out = 8'h2F;
                    16'h1E12: data_out = 8'h30;
                    16'h1E13: data_out = 8'h31;
                    16'h1E14: data_out = 8'h32;
                    16'h1E15: data_out = 8'h33;
                    16'h1E16: data_out = 8'h34;
                    16'h1E17: data_out = 8'h35;
                    16'h1E18: data_out = 8'h36;
                    16'h1E19: data_out = 8'h37;
                    16'h1E1A: data_out = 8'h38;
                    16'h1E1B: data_out = 8'h39;
                    16'h1E1C: data_out = 8'h3A;
                    16'h1E1D: data_out = 8'h3B;
                    16'h1E1E: data_out = 8'h3C;
                    16'h1E1F: data_out = 8'h3D;
                    16'h1E20: data_out = 8'h3E;
                    16'h1E21: data_out = 8'h3F;
                    16'h1E22: data_out = 8'h40;
                    16'h1E23: data_out = 8'h41;
                    16'h1E24: data_out = 8'h42;
                    16'h1E25: data_out = 8'h43;
                    16'h1E26: data_out = 8'h44;
                    16'h1E27: data_out = 8'h45;
                    16'h1E28: data_out = 8'h46;
                    16'h1E29: data_out = 8'h47;
                    16'h1E2A: data_out = 8'h48;
                    16'h1E2B: data_out = 8'h49;
                    16'h1E2C: data_out = 8'h4A;
                    16'h1E2D: data_out = 8'h4B;
                    16'h1E2E: data_out = 8'h4C;
                    16'h1E2F: data_out = 8'h4D;
                    16'h1E30: data_out = 8'h4E;
                    16'h1E31: data_out = 8'h4F;
                    16'h1E32: data_out = 8'h50;
                    16'h1E33: data_out = 8'h51;
                    16'h1E34: data_out = 8'h52;
                    16'h1E35: data_out = 8'h53;
                    16'h1E36: data_out = 8'h54;
                    16'h1E37: data_out = 8'h55;
                    16'h1E38: data_out = 8'h56;
                    16'h1E39: data_out = 8'h57;
                    16'h1E3A: data_out = 8'h58;
                    16'h1E3B: data_out = 8'h59;
                    16'h1E3C: data_out = 8'h5A;
                    16'h1E3D: data_out = 8'h5B;
                    16'h1E3E: data_out = 8'h5C;
                    16'h1E3F: data_out = 8'h5D;
                    16'h1E40: data_out = 8'h5E;
                    16'h1E41: data_out = 8'h5F;
                    16'h1E42: data_out = 8'h60;
                    16'h1E43: data_out = 8'h61;
                    16'h1E44: data_out = 8'h62;
                    16'h1E45: data_out = 8'h63;
                    16'h1E46: data_out = 8'h64;
                    16'h1E47: data_out = 8'h65;
                    16'h1E48: data_out = 8'h66;
                    16'h1E49: data_out = 8'h67;
                    16'h1E4A: data_out = 8'h68;
                    16'h1E4B: data_out = 8'h69;
                    16'h1E4C: data_out = 8'h6A;
                    16'h1E4D: data_out = 8'h6B;
                    16'h1E4E: data_out = 8'h6C;
                    16'h1E4F: data_out = 8'h6D;
                    16'h1E50: data_out = 8'h6E;
                    16'h1E51: data_out = 8'h6F;
                    16'h1E52: data_out = 8'h70;
                    16'h1E53: data_out = 8'h71;
                    16'h1E54: data_out = 8'h72;
                    16'h1E55: data_out = 8'h73;
                    16'h1E56: data_out = 8'h74;
                    16'h1E57: data_out = 8'h75;
                    16'h1E58: data_out = 8'h76;
                    16'h1E59: data_out = 8'h77;
                    16'h1E5A: data_out = 8'h78;
                    16'h1E5B: data_out = 8'h79;
                    16'h1E5C: data_out = 8'h7A;
                    16'h1E5D: data_out = 8'h7B;
                    16'h1E5E: data_out = 8'h7C;
                    16'h1E5F: data_out = 8'h7D;
                    16'h1E60: data_out = 8'h7E;
                    16'h1E61: data_out = 8'h7F;
                    16'h1E62: data_out = 8'h80;
                    16'h1E63: data_out = 8'h81;
                    16'h1E64: data_out = 8'h82;
                    16'h1E65: data_out = 8'h83;
                    16'h1E66: data_out = 8'h84;
                    16'h1E67: data_out = 8'h85;
                    16'h1E68: data_out = 8'h86;
                    16'h1E69: data_out = 8'h87;
                    16'h1E6A: data_out = 8'h88;
                    16'h1E6B: data_out = 8'h89;
                    16'h1E6C: data_out = 8'h8A;
                    16'h1E6D: data_out = 8'h8B;
                    16'h1E6E: data_out = 8'h8C;
                    16'h1E6F: data_out = 8'h8D;
                    16'h1E70: data_out = 8'h8E;
                    16'h1E71: data_out = 8'h8F;
                    16'h1E72: data_out = 8'h90;
                    16'h1E73: data_out = 8'h91;
                    16'h1E74: data_out = 8'h92;
                    16'h1E75: data_out = 8'h93;
                    16'h1E76: data_out = 8'h94;
                    16'h1E77: data_out = 8'h95;
                    16'h1E78: data_out = 8'h96;
                    16'h1E79: data_out = 8'h97;
                    16'h1E7A: data_out = 8'h98;
                    16'h1E7B: data_out = 8'h99;
                    16'h1E7C: data_out = 8'h9A;
                    16'h1E7D: data_out = 8'h9B;
                    16'h1E7E: data_out = 8'h9C;
                    16'h1E7F: data_out = 8'h9D;
                    16'h1E80: data_out = 8'h1E;
                    16'h1E81: data_out = 8'h1D;
                    16'h1E82: data_out = 8'h1C;
                    16'h1E83: data_out = 8'h1B;
                    16'h1E84: data_out = 8'h1A;
                    16'h1E85: data_out = 8'h19;
                    16'h1E86: data_out = 8'h18;
                    16'h1E87: data_out = 8'h17;
                    16'h1E88: data_out = 8'h16;
                    16'h1E89: data_out = 8'h15;
                    16'h1E8A: data_out = 8'h14;
                    16'h1E8B: data_out = 8'h13;
                    16'h1E8C: data_out = 8'h12;
                    16'h1E8D: data_out = 8'h11;
                    16'h1E8E: data_out = 8'h10;
                    16'h1E8F: data_out = 8'hF;
                    16'h1E90: data_out = 8'hE;
                    16'h1E91: data_out = 8'hD;
                    16'h1E92: data_out = 8'hC;
                    16'h1E93: data_out = 8'hB;
                    16'h1E94: data_out = 8'hA;
                    16'h1E95: data_out = 8'h9;
                    16'h1E96: data_out = 8'h8;
                    16'h1E97: data_out = 8'h7;
                    16'h1E98: data_out = 8'h6;
                    16'h1E99: data_out = 8'h5;
                    16'h1E9A: data_out = 8'h4;
                    16'h1E9B: data_out = 8'h3;
                    16'h1E9C: data_out = 8'h2;
                    16'h1E9D: data_out = 8'h1;
                    16'h1E9E: data_out = 8'h0;
                    16'h1E9F: data_out = 8'h81;
                    16'h1EA0: data_out = 8'h82;
                    16'h1EA1: data_out = 8'h83;
                    16'h1EA2: data_out = 8'h84;
                    16'h1EA3: data_out = 8'h85;
                    16'h1EA4: data_out = 8'h86;
                    16'h1EA5: data_out = 8'h87;
                    16'h1EA6: data_out = 8'h88;
                    16'h1EA7: data_out = 8'h89;
                    16'h1EA8: data_out = 8'h8A;
                    16'h1EA9: data_out = 8'h8B;
                    16'h1EAA: data_out = 8'h8C;
                    16'h1EAB: data_out = 8'h8D;
                    16'h1EAC: data_out = 8'h8E;
                    16'h1EAD: data_out = 8'h8F;
                    16'h1EAE: data_out = 8'h90;
                    16'h1EAF: data_out = 8'h91;
                    16'h1EB0: data_out = 8'h92;
                    16'h1EB1: data_out = 8'h93;
                    16'h1EB2: data_out = 8'h94;
                    16'h1EB3: data_out = 8'h95;
                    16'h1EB4: data_out = 8'h96;
                    16'h1EB5: data_out = 8'h97;
                    16'h1EB6: data_out = 8'h98;
                    16'h1EB7: data_out = 8'h99;
                    16'h1EB8: data_out = 8'h9A;
                    16'h1EB9: data_out = 8'h9B;
                    16'h1EBA: data_out = 8'h9C;
                    16'h1EBB: data_out = 8'h9D;
                    16'h1EBC: data_out = 8'h9E;
                    16'h1EBD: data_out = 8'h9F;
                    16'h1EBE: data_out = 8'hA0;
                    16'h1EBF: data_out = 8'hA1;
                    16'h1EC0: data_out = 8'hA2;
                    16'h1EC1: data_out = 8'hA3;
                    16'h1EC2: data_out = 8'hA4;
                    16'h1EC3: data_out = 8'hA5;
                    16'h1EC4: data_out = 8'hA6;
                    16'h1EC5: data_out = 8'hA7;
                    16'h1EC6: data_out = 8'hA8;
                    16'h1EC7: data_out = 8'hA9;
                    16'h1EC8: data_out = 8'hAA;
                    16'h1EC9: data_out = 8'hAB;
                    16'h1ECA: data_out = 8'hAC;
                    16'h1ECB: data_out = 8'hAD;
                    16'h1ECC: data_out = 8'hAE;
                    16'h1ECD: data_out = 8'hAF;
                    16'h1ECE: data_out = 8'hB0;
                    16'h1ECF: data_out = 8'hB1;
                    16'h1ED0: data_out = 8'hB2;
                    16'h1ED1: data_out = 8'hB3;
                    16'h1ED2: data_out = 8'hB4;
                    16'h1ED3: data_out = 8'hB5;
                    16'h1ED4: data_out = 8'hB6;
                    16'h1ED5: data_out = 8'hB7;
                    16'h1ED6: data_out = 8'hB8;
                    16'h1ED7: data_out = 8'hB9;
                    16'h1ED8: data_out = 8'hBA;
                    16'h1ED9: data_out = 8'hBB;
                    16'h1EDA: data_out = 8'hBC;
                    16'h1EDB: data_out = 8'hBD;
                    16'h1EDC: data_out = 8'hBE;
                    16'h1EDD: data_out = 8'hBF;
                    16'h1EDE: data_out = 8'hC0;
                    16'h1EDF: data_out = 8'hC1;
                    16'h1EE0: data_out = 8'hC2;
                    16'h1EE1: data_out = 8'hC3;
                    16'h1EE2: data_out = 8'hC4;
                    16'h1EE3: data_out = 8'hC5;
                    16'h1EE4: data_out = 8'hC6;
                    16'h1EE5: data_out = 8'hC7;
                    16'h1EE6: data_out = 8'hC8;
                    16'h1EE7: data_out = 8'hC9;
                    16'h1EE8: data_out = 8'hCA;
                    16'h1EE9: data_out = 8'hCB;
                    16'h1EEA: data_out = 8'hCC;
                    16'h1EEB: data_out = 8'hCD;
                    16'h1EEC: data_out = 8'hCE;
                    16'h1EED: data_out = 8'hCF;
                    16'h1EEE: data_out = 8'hD0;
                    16'h1EEF: data_out = 8'hD1;
                    16'h1EF0: data_out = 8'hD2;
                    16'h1EF1: data_out = 8'hD3;
                    16'h1EF2: data_out = 8'hD4;
                    16'h1EF3: data_out = 8'hD5;
                    16'h1EF4: data_out = 8'hD6;
                    16'h1EF5: data_out = 8'hD7;
                    16'h1EF6: data_out = 8'hD8;
                    16'h1EF7: data_out = 8'hD9;
                    16'h1EF8: data_out = 8'hDA;
                    16'h1EF9: data_out = 8'hDB;
                    16'h1EFA: data_out = 8'hDC;
                    16'h1EFB: data_out = 8'hDD;
                    16'h1EFC: data_out = 8'hDE;
                    16'h1EFD: data_out = 8'hDF;
                    16'h1EFE: data_out = 8'hE0;
                    16'h1EFF: data_out = 8'hE1;
                    16'h1F00: data_out = 8'h1F;
                    16'h1F01: data_out = 8'h20;
                    16'h1F02: data_out = 8'h21;
                    16'h1F03: data_out = 8'h22;
                    16'h1F04: data_out = 8'h23;
                    16'h1F05: data_out = 8'h24;
                    16'h1F06: data_out = 8'h25;
                    16'h1F07: data_out = 8'h26;
                    16'h1F08: data_out = 8'h27;
                    16'h1F09: data_out = 8'h28;
                    16'h1F0A: data_out = 8'h29;
                    16'h1F0B: data_out = 8'h2A;
                    16'h1F0C: data_out = 8'h2B;
                    16'h1F0D: data_out = 8'h2C;
                    16'h1F0E: data_out = 8'h2D;
                    16'h1F0F: data_out = 8'h2E;
                    16'h1F10: data_out = 8'h2F;
                    16'h1F11: data_out = 8'h30;
                    16'h1F12: data_out = 8'h31;
                    16'h1F13: data_out = 8'h32;
                    16'h1F14: data_out = 8'h33;
                    16'h1F15: data_out = 8'h34;
                    16'h1F16: data_out = 8'h35;
                    16'h1F17: data_out = 8'h36;
                    16'h1F18: data_out = 8'h37;
                    16'h1F19: data_out = 8'h38;
                    16'h1F1A: data_out = 8'h39;
                    16'h1F1B: data_out = 8'h3A;
                    16'h1F1C: data_out = 8'h3B;
                    16'h1F1D: data_out = 8'h3C;
                    16'h1F1E: data_out = 8'h3D;
                    16'h1F1F: data_out = 8'h3E;
                    16'h1F20: data_out = 8'h3F;
                    16'h1F21: data_out = 8'h40;
                    16'h1F22: data_out = 8'h41;
                    16'h1F23: data_out = 8'h42;
                    16'h1F24: data_out = 8'h43;
                    16'h1F25: data_out = 8'h44;
                    16'h1F26: data_out = 8'h45;
                    16'h1F27: data_out = 8'h46;
                    16'h1F28: data_out = 8'h47;
                    16'h1F29: data_out = 8'h48;
                    16'h1F2A: data_out = 8'h49;
                    16'h1F2B: data_out = 8'h4A;
                    16'h1F2C: data_out = 8'h4B;
                    16'h1F2D: data_out = 8'h4C;
                    16'h1F2E: data_out = 8'h4D;
                    16'h1F2F: data_out = 8'h4E;
                    16'h1F30: data_out = 8'h4F;
                    16'h1F31: data_out = 8'h50;
                    16'h1F32: data_out = 8'h51;
                    16'h1F33: data_out = 8'h52;
                    16'h1F34: data_out = 8'h53;
                    16'h1F35: data_out = 8'h54;
                    16'h1F36: data_out = 8'h55;
                    16'h1F37: data_out = 8'h56;
                    16'h1F38: data_out = 8'h57;
                    16'h1F39: data_out = 8'h58;
                    16'h1F3A: data_out = 8'h59;
                    16'h1F3B: data_out = 8'h5A;
                    16'h1F3C: data_out = 8'h5B;
                    16'h1F3D: data_out = 8'h5C;
                    16'h1F3E: data_out = 8'h5D;
                    16'h1F3F: data_out = 8'h5E;
                    16'h1F40: data_out = 8'h5F;
                    16'h1F41: data_out = 8'h60;
                    16'h1F42: data_out = 8'h61;
                    16'h1F43: data_out = 8'h62;
                    16'h1F44: data_out = 8'h63;
                    16'h1F45: data_out = 8'h64;
                    16'h1F46: data_out = 8'h65;
                    16'h1F47: data_out = 8'h66;
                    16'h1F48: data_out = 8'h67;
                    16'h1F49: data_out = 8'h68;
                    16'h1F4A: data_out = 8'h69;
                    16'h1F4B: data_out = 8'h6A;
                    16'h1F4C: data_out = 8'h6B;
                    16'h1F4D: data_out = 8'h6C;
                    16'h1F4E: data_out = 8'h6D;
                    16'h1F4F: data_out = 8'h6E;
                    16'h1F50: data_out = 8'h6F;
                    16'h1F51: data_out = 8'h70;
                    16'h1F52: data_out = 8'h71;
                    16'h1F53: data_out = 8'h72;
                    16'h1F54: data_out = 8'h73;
                    16'h1F55: data_out = 8'h74;
                    16'h1F56: data_out = 8'h75;
                    16'h1F57: data_out = 8'h76;
                    16'h1F58: data_out = 8'h77;
                    16'h1F59: data_out = 8'h78;
                    16'h1F5A: data_out = 8'h79;
                    16'h1F5B: data_out = 8'h7A;
                    16'h1F5C: data_out = 8'h7B;
                    16'h1F5D: data_out = 8'h7C;
                    16'h1F5E: data_out = 8'h7D;
                    16'h1F5F: data_out = 8'h7E;
                    16'h1F60: data_out = 8'h7F;
                    16'h1F61: data_out = 8'h80;
                    16'h1F62: data_out = 8'h81;
                    16'h1F63: data_out = 8'h82;
                    16'h1F64: data_out = 8'h83;
                    16'h1F65: data_out = 8'h84;
                    16'h1F66: data_out = 8'h85;
                    16'h1F67: data_out = 8'h86;
                    16'h1F68: data_out = 8'h87;
                    16'h1F69: data_out = 8'h88;
                    16'h1F6A: data_out = 8'h89;
                    16'h1F6B: data_out = 8'h8A;
                    16'h1F6C: data_out = 8'h8B;
                    16'h1F6D: data_out = 8'h8C;
                    16'h1F6E: data_out = 8'h8D;
                    16'h1F6F: data_out = 8'h8E;
                    16'h1F70: data_out = 8'h8F;
                    16'h1F71: data_out = 8'h90;
                    16'h1F72: data_out = 8'h91;
                    16'h1F73: data_out = 8'h92;
                    16'h1F74: data_out = 8'h93;
                    16'h1F75: data_out = 8'h94;
                    16'h1F76: data_out = 8'h95;
                    16'h1F77: data_out = 8'h96;
                    16'h1F78: data_out = 8'h97;
                    16'h1F79: data_out = 8'h98;
                    16'h1F7A: data_out = 8'h99;
                    16'h1F7B: data_out = 8'h9A;
                    16'h1F7C: data_out = 8'h9B;
                    16'h1F7D: data_out = 8'h9C;
                    16'h1F7E: data_out = 8'h9D;
                    16'h1F7F: data_out = 8'h9E;
                    16'h1F80: data_out = 8'h1F;
                    16'h1F81: data_out = 8'h1E;
                    16'h1F82: data_out = 8'h1D;
                    16'h1F83: data_out = 8'h1C;
                    16'h1F84: data_out = 8'h1B;
                    16'h1F85: data_out = 8'h1A;
                    16'h1F86: data_out = 8'h19;
                    16'h1F87: data_out = 8'h18;
                    16'h1F88: data_out = 8'h17;
                    16'h1F89: data_out = 8'h16;
                    16'h1F8A: data_out = 8'h15;
                    16'h1F8B: data_out = 8'h14;
                    16'h1F8C: data_out = 8'h13;
                    16'h1F8D: data_out = 8'h12;
                    16'h1F8E: data_out = 8'h11;
                    16'h1F8F: data_out = 8'h10;
                    16'h1F90: data_out = 8'hF;
                    16'h1F91: data_out = 8'hE;
                    16'h1F92: data_out = 8'hD;
                    16'h1F93: data_out = 8'hC;
                    16'h1F94: data_out = 8'hB;
                    16'h1F95: data_out = 8'hA;
                    16'h1F96: data_out = 8'h9;
                    16'h1F97: data_out = 8'h8;
                    16'h1F98: data_out = 8'h7;
                    16'h1F99: data_out = 8'h6;
                    16'h1F9A: data_out = 8'h5;
                    16'h1F9B: data_out = 8'h4;
                    16'h1F9C: data_out = 8'h3;
                    16'h1F9D: data_out = 8'h2;
                    16'h1F9E: data_out = 8'h1;
                    16'h1F9F: data_out = 8'h0;
                    16'h1FA0: data_out = 8'h81;
                    16'h1FA1: data_out = 8'h82;
                    16'h1FA2: data_out = 8'h83;
                    16'h1FA3: data_out = 8'h84;
                    16'h1FA4: data_out = 8'h85;
                    16'h1FA5: data_out = 8'h86;
                    16'h1FA6: data_out = 8'h87;
                    16'h1FA7: data_out = 8'h88;
                    16'h1FA8: data_out = 8'h89;
                    16'h1FA9: data_out = 8'h8A;
                    16'h1FAA: data_out = 8'h8B;
                    16'h1FAB: data_out = 8'h8C;
                    16'h1FAC: data_out = 8'h8D;
                    16'h1FAD: data_out = 8'h8E;
                    16'h1FAE: data_out = 8'h8F;
                    16'h1FAF: data_out = 8'h90;
                    16'h1FB0: data_out = 8'h91;
                    16'h1FB1: data_out = 8'h92;
                    16'h1FB2: data_out = 8'h93;
                    16'h1FB3: data_out = 8'h94;
                    16'h1FB4: data_out = 8'h95;
                    16'h1FB5: data_out = 8'h96;
                    16'h1FB6: data_out = 8'h97;
                    16'h1FB7: data_out = 8'h98;
                    16'h1FB8: data_out = 8'h99;
                    16'h1FB9: data_out = 8'h9A;
                    16'h1FBA: data_out = 8'h9B;
                    16'h1FBB: data_out = 8'h9C;
                    16'h1FBC: data_out = 8'h9D;
                    16'h1FBD: data_out = 8'h9E;
                    16'h1FBE: data_out = 8'h9F;
                    16'h1FBF: data_out = 8'hA0;
                    16'h1FC0: data_out = 8'hA1;
                    16'h1FC1: data_out = 8'hA2;
                    16'h1FC2: data_out = 8'hA3;
                    16'h1FC3: data_out = 8'hA4;
                    16'h1FC4: data_out = 8'hA5;
                    16'h1FC5: data_out = 8'hA6;
                    16'h1FC6: data_out = 8'hA7;
                    16'h1FC7: data_out = 8'hA8;
                    16'h1FC8: data_out = 8'hA9;
                    16'h1FC9: data_out = 8'hAA;
                    16'h1FCA: data_out = 8'hAB;
                    16'h1FCB: data_out = 8'hAC;
                    16'h1FCC: data_out = 8'hAD;
                    16'h1FCD: data_out = 8'hAE;
                    16'h1FCE: data_out = 8'hAF;
                    16'h1FCF: data_out = 8'hB0;
                    16'h1FD0: data_out = 8'hB1;
                    16'h1FD1: data_out = 8'hB2;
                    16'h1FD2: data_out = 8'hB3;
                    16'h1FD3: data_out = 8'hB4;
                    16'h1FD4: data_out = 8'hB5;
                    16'h1FD5: data_out = 8'hB6;
                    16'h1FD6: data_out = 8'hB7;
                    16'h1FD7: data_out = 8'hB8;
                    16'h1FD8: data_out = 8'hB9;
                    16'h1FD9: data_out = 8'hBA;
                    16'h1FDA: data_out = 8'hBB;
                    16'h1FDB: data_out = 8'hBC;
                    16'h1FDC: data_out = 8'hBD;
                    16'h1FDD: data_out = 8'hBE;
                    16'h1FDE: data_out = 8'hBF;
                    16'h1FDF: data_out = 8'hC0;
                    16'h1FE0: data_out = 8'hC1;
                    16'h1FE1: data_out = 8'hC2;
                    16'h1FE2: data_out = 8'hC3;
                    16'h1FE3: data_out = 8'hC4;
                    16'h1FE4: data_out = 8'hC5;
                    16'h1FE5: data_out = 8'hC6;
                    16'h1FE6: data_out = 8'hC7;
                    16'h1FE7: data_out = 8'hC8;
                    16'h1FE8: data_out = 8'hC9;
                    16'h1FE9: data_out = 8'hCA;
                    16'h1FEA: data_out = 8'hCB;
                    16'h1FEB: data_out = 8'hCC;
                    16'h1FEC: data_out = 8'hCD;
                    16'h1FED: data_out = 8'hCE;
                    16'h1FEE: data_out = 8'hCF;
                    16'h1FEF: data_out = 8'hD0;
                    16'h1FF0: data_out = 8'hD1;
                    16'h1FF1: data_out = 8'hD2;
                    16'h1FF2: data_out = 8'hD3;
                    16'h1FF3: data_out = 8'hD4;
                    16'h1FF4: data_out = 8'hD5;
                    16'h1FF5: data_out = 8'hD6;
                    16'h1FF6: data_out = 8'hD7;
                    16'h1FF7: data_out = 8'hD8;
                    16'h1FF8: data_out = 8'hD9;
                    16'h1FF9: data_out = 8'hDA;
                    16'h1FFA: data_out = 8'hDB;
                    16'h1FFB: data_out = 8'hDC;
                    16'h1FFC: data_out = 8'hDD;
                    16'h1FFD: data_out = 8'hDE;
                    16'h1FFE: data_out = 8'hDF;
                    16'h1FFF: data_out = 8'hE0;
                    16'h2000: data_out = 8'h20;
                    16'h2001: data_out = 8'h21;
                    16'h2002: data_out = 8'h22;
                    16'h2003: data_out = 8'h23;
                    16'h2004: data_out = 8'h24;
                    16'h2005: data_out = 8'h25;
                    16'h2006: data_out = 8'h26;
                    16'h2007: data_out = 8'h27;
                    16'h2008: data_out = 8'h28;
                    16'h2009: data_out = 8'h29;
                    16'h200A: data_out = 8'h2A;
                    16'h200B: data_out = 8'h2B;
                    16'h200C: data_out = 8'h2C;
                    16'h200D: data_out = 8'h2D;
                    16'h200E: data_out = 8'h2E;
                    16'h200F: data_out = 8'h2F;
                    16'h2010: data_out = 8'h30;
                    16'h2011: data_out = 8'h31;
                    16'h2012: data_out = 8'h32;
                    16'h2013: data_out = 8'h33;
                    16'h2014: data_out = 8'h34;
                    16'h2015: data_out = 8'h35;
                    16'h2016: data_out = 8'h36;
                    16'h2017: data_out = 8'h37;
                    16'h2018: data_out = 8'h38;
                    16'h2019: data_out = 8'h39;
                    16'h201A: data_out = 8'h3A;
                    16'h201B: data_out = 8'h3B;
                    16'h201C: data_out = 8'h3C;
                    16'h201D: data_out = 8'h3D;
                    16'h201E: data_out = 8'h3E;
                    16'h201F: data_out = 8'h3F;
                    16'h2020: data_out = 8'h40;
                    16'h2021: data_out = 8'h41;
                    16'h2022: data_out = 8'h42;
                    16'h2023: data_out = 8'h43;
                    16'h2024: data_out = 8'h44;
                    16'h2025: data_out = 8'h45;
                    16'h2026: data_out = 8'h46;
                    16'h2027: data_out = 8'h47;
                    16'h2028: data_out = 8'h48;
                    16'h2029: data_out = 8'h49;
                    16'h202A: data_out = 8'h4A;
                    16'h202B: data_out = 8'h4B;
                    16'h202C: data_out = 8'h4C;
                    16'h202D: data_out = 8'h4D;
                    16'h202E: data_out = 8'h4E;
                    16'h202F: data_out = 8'h4F;
                    16'h2030: data_out = 8'h50;
                    16'h2031: data_out = 8'h51;
                    16'h2032: data_out = 8'h52;
                    16'h2033: data_out = 8'h53;
                    16'h2034: data_out = 8'h54;
                    16'h2035: data_out = 8'h55;
                    16'h2036: data_out = 8'h56;
                    16'h2037: data_out = 8'h57;
                    16'h2038: data_out = 8'h58;
                    16'h2039: data_out = 8'h59;
                    16'h203A: data_out = 8'h5A;
                    16'h203B: data_out = 8'h5B;
                    16'h203C: data_out = 8'h5C;
                    16'h203D: data_out = 8'h5D;
                    16'h203E: data_out = 8'h5E;
                    16'h203F: data_out = 8'h5F;
                    16'h2040: data_out = 8'h60;
                    16'h2041: data_out = 8'h61;
                    16'h2042: data_out = 8'h62;
                    16'h2043: data_out = 8'h63;
                    16'h2044: data_out = 8'h64;
                    16'h2045: data_out = 8'h65;
                    16'h2046: data_out = 8'h66;
                    16'h2047: data_out = 8'h67;
                    16'h2048: data_out = 8'h68;
                    16'h2049: data_out = 8'h69;
                    16'h204A: data_out = 8'h6A;
                    16'h204B: data_out = 8'h6B;
                    16'h204C: data_out = 8'h6C;
                    16'h204D: data_out = 8'h6D;
                    16'h204E: data_out = 8'h6E;
                    16'h204F: data_out = 8'h6F;
                    16'h2050: data_out = 8'h70;
                    16'h2051: data_out = 8'h71;
                    16'h2052: data_out = 8'h72;
                    16'h2053: data_out = 8'h73;
                    16'h2054: data_out = 8'h74;
                    16'h2055: data_out = 8'h75;
                    16'h2056: data_out = 8'h76;
                    16'h2057: data_out = 8'h77;
                    16'h2058: data_out = 8'h78;
                    16'h2059: data_out = 8'h79;
                    16'h205A: data_out = 8'h7A;
                    16'h205B: data_out = 8'h7B;
                    16'h205C: data_out = 8'h7C;
                    16'h205D: data_out = 8'h7D;
                    16'h205E: data_out = 8'h7E;
                    16'h205F: data_out = 8'h7F;
                    16'h2060: data_out = 8'h80;
                    16'h2061: data_out = 8'h81;
                    16'h2062: data_out = 8'h82;
                    16'h2063: data_out = 8'h83;
                    16'h2064: data_out = 8'h84;
                    16'h2065: data_out = 8'h85;
                    16'h2066: data_out = 8'h86;
                    16'h2067: data_out = 8'h87;
                    16'h2068: data_out = 8'h88;
                    16'h2069: data_out = 8'h89;
                    16'h206A: data_out = 8'h8A;
                    16'h206B: data_out = 8'h8B;
                    16'h206C: data_out = 8'h8C;
                    16'h206D: data_out = 8'h8D;
                    16'h206E: data_out = 8'h8E;
                    16'h206F: data_out = 8'h8F;
                    16'h2070: data_out = 8'h90;
                    16'h2071: data_out = 8'h91;
                    16'h2072: data_out = 8'h92;
                    16'h2073: data_out = 8'h93;
                    16'h2074: data_out = 8'h94;
                    16'h2075: data_out = 8'h95;
                    16'h2076: data_out = 8'h96;
                    16'h2077: data_out = 8'h97;
                    16'h2078: data_out = 8'h98;
                    16'h2079: data_out = 8'h99;
                    16'h207A: data_out = 8'h9A;
                    16'h207B: data_out = 8'h9B;
                    16'h207C: data_out = 8'h9C;
                    16'h207D: data_out = 8'h9D;
                    16'h207E: data_out = 8'h9E;
                    16'h207F: data_out = 8'h9F;
                    16'h2080: data_out = 8'h20;
                    16'h2081: data_out = 8'h1F;
                    16'h2082: data_out = 8'h1E;
                    16'h2083: data_out = 8'h1D;
                    16'h2084: data_out = 8'h1C;
                    16'h2085: data_out = 8'h1B;
                    16'h2086: data_out = 8'h1A;
                    16'h2087: data_out = 8'h19;
                    16'h2088: data_out = 8'h18;
                    16'h2089: data_out = 8'h17;
                    16'h208A: data_out = 8'h16;
                    16'h208B: data_out = 8'h15;
                    16'h208C: data_out = 8'h14;
                    16'h208D: data_out = 8'h13;
                    16'h208E: data_out = 8'h12;
                    16'h208F: data_out = 8'h11;
                    16'h2090: data_out = 8'h10;
                    16'h2091: data_out = 8'hF;
                    16'h2092: data_out = 8'hE;
                    16'h2093: data_out = 8'hD;
                    16'h2094: data_out = 8'hC;
                    16'h2095: data_out = 8'hB;
                    16'h2096: data_out = 8'hA;
                    16'h2097: data_out = 8'h9;
                    16'h2098: data_out = 8'h8;
                    16'h2099: data_out = 8'h7;
                    16'h209A: data_out = 8'h6;
                    16'h209B: data_out = 8'h5;
                    16'h209C: data_out = 8'h4;
                    16'h209D: data_out = 8'h3;
                    16'h209E: data_out = 8'h2;
                    16'h209F: data_out = 8'h1;
                    16'h20A0: data_out = 8'h0;
                    16'h20A1: data_out = 8'h81;
                    16'h20A2: data_out = 8'h82;
                    16'h20A3: data_out = 8'h83;
                    16'h20A4: data_out = 8'h84;
                    16'h20A5: data_out = 8'h85;
                    16'h20A6: data_out = 8'h86;
                    16'h20A7: data_out = 8'h87;
                    16'h20A8: data_out = 8'h88;
                    16'h20A9: data_out = 8'h89;
                    16'h20AA: data_out = 8'h8A;
                    16'h20AB: data_out = 8'h8B;
                    16'h20AC: data_out = 8'h8C;
                    16'h20AD: data_out = 8'h8D;
                    16'h20AE: data_out = 8'h8E;
                    16'h20AF: data_out = 8'h8F;
                    16'h20B0: data_out = 8'h90;
                    16'h20B1: data_out = 8'h91;
                    16'h20B2: data_out = 8'h92;
                    16'h20B3: data_out = 8'h93;
                    16'h20B4: data_out = 8'h94;
                    16'h20B5: data_out = 8'h95;
                    16'h20B6: data_out = 8'h96;
                    16'h20B7: data_out = 8'h97;
                    16'h20B8: data_out = 8'h98;
                    16'h20B9: data_out = 8'h99;
                    16'h20BA: data_out = 8'h9A;
                    16'h20BB: data_out = 8'h9B;
                    16'h20BC: data_out = 8'h9C;
                    16'h20BD: data_out = 8'h9D;
                    16'h20BE: data_out = 8'h9E;
                    16'h20BF: data_out = 8'h9F;
                    16'h20C0: data_out = 8'hA0;
                    16'h20C1: data_out = 8'hA1;
                    16'h20C2: data_out = 8'hA2;
                    16'h20C3: data_out = 8'hA3;
                    16'h20C4: data_out = 8'hA4;
                    16'h20C5: data_out = 8'hA5;
                    16'h20C6: data_out = 8'hA6;
                    16'h20C7: data_out = 8'hA7;
                    16'h20C8: data_out = 8'hA8;
                    16'h20C9: data_out = 8'hA9;
                    16'h20CA: data_out = 8'hAA;
                    16'h20CB: data_out = 8'hAB;
                    16'h20CC: data_out = 8'hAC;
                    16'h20CD: data_out = 8'hAD;
                    16'h20CE: data_out = 8'hAE;
                    16'h20CF: data_out = 8'hAF;
                    16'h20D0: data_out = 8'hB0;
                    16'h20D1: data_out = 8'hB1;
                    16'h20D2: data_out = 8'hB2;
                    16'h20D3: data_out = 8'hB3;
                    16'h20D4: data_out = 8'hB4;
                    16'h20D5: data_out = 8'hB5;
                    16'h20D6: data_out = 8'hB6;
                    16'h20D7: data_out = 8'hB7;
                    16'h20D8: data_out = 8'hB8;
                    16'h20D9: data_out = 8'hB9;
                    16'h20DA: data_out = 8'hBA;
                    16'h20DB: data_out = 8'hBB;
                    16'h20DC: data_out = 8'hBC;
                    16'h20DD: data_out = 8'hBD;
                    16'h20DE: data_out = 8'hBE;
                    16'h20DF: data_out = 8'hBF;
                    16'h20E0: data_out = 8'hC0;
                    16'h20E1: data_out = 8'hC1;
                    16'h20E2: data_out = 8'hC2;
                    16'h20E3: data_out = 8'hC3;
                    16'h20E4: data_out = 8'hC4;
                    16'h20E5: data_out = 8'hC5;
                    16'h20E6: data_out = 8'hC6;
                    16'h20E7: data_out = 8'hC7;
                    16'h20E8: data_out = 8'hC8;
                    16'h20E9: data_out = 8'hC9;
                    16'h20EA: data_out = 8'hCA;
                    16'h20EB: data_out = 8'hCB;
                    16'h20EC: data_out = 8'hCC;
                    16'h20ED: data_out = 8'hCD;
                    16'h20EE: data_out = 8'hCE;
                    16'h20EF: data_out = 8'hCF;
                    16'h20F0: data_out = 8'hD0;
                    16'h20F1: data_out = 8'hD1;
                    16'h20F2: data_out = 8'hD2;
                    16'h20F3: data_out = 8'hD3;
                    16'h20F4: data_out = 8'hD4;
                    16'h20F5: data_out = 8'hD5;
                    16'h20F6: data_out = 8'hD6;
                    16'h20F7: data_out = 8'hD7;
                    16'h20F8: data_out = 8'hD8;
                    16'h20F9: data_out = 8'hD9;
                    16'h20FA: data_out = 8'hDA;
                    16'h20FB: data_out = 8'hDB;
                    16'h20FC: data_out = 8'hDC;
                    16'h20FD: data_out = 8'hDD;
                    16'h20FE: data_out = 8'hDE;
                    16'h20FF: data_out = 8'hDF;
                    16'h2100: data_out = 8'h21;
                    16'h2101: data_out = 8'h22;
                    16'h2102: data_out = 8'h23;
                    16'h2103: data_out = 8'h24;
                    16'h2104: data_out = 8'h25;
                    16'h2105: data_out = 8'h26;
                    16'h2106: data_out = 8'h27;
                    16'h2107: data_out = 8'h28;
                    16'h2108: data_out = 8'h29;
                    16'h2109: data_out = 8'h2A;
                    16'h210A: data_out = 8'h2B;
                    16'h210B: data_out = 8'h2C;
                    16'h210C: data_out = 8'h2D;
                    16'h210D: data_out = 8'h2E;
                    16'h210E: data_out = 8'h2F;
                    16'h210F: data_out = 8'h30;
                    16'h2110: data_out = 8'h31;
                    16'h2111: data_out = 8'h32;
                    16'h2112: data_out = 8'h33;
                    16'h2113: data_out = 8'h34;
                    16'h2114: data_out = 8'h35;
                    16'h2115: data_out = 8'h36;
                    16'h2116: data_out = 8'h37;
                    16'h2117: data_out = 8'h38;
                    16'h2118: data_out = 8'h39;
                    16'h2119: data_out = 8'h3A;
                    16'h211A: data_out = 8'h3B;
                    16'h211B: data_out = 8'h3C;
                    16'h211C: data_out = 8'h3D;
                    16'h211D: data_out = 8'h3E;
                    16'h211E: data_out = 8'h3F;
                    16'h211F: data_out = 8'h40;
                    16'h2120: data_out = 8'h41;
                    16'h2121: data_out = 8'h42;
                    16'h2122: data_out = 8'h43;
                    16'h2123: data_out = 8'h44;
                    16'h2124: data_out = 8'h45;
                    16'h2125: data_out = 8'h46;
                    16'h2126: data_out = 8'h47;
                    16'h2127: data_out = 8'h48;
                    16'h2128: data_out = 8'h49;
                    16'h2129: data_out = 8'h4A;
                    16'h212A: data_out = 8'h4B;
                    16'h212B: data_out = 8'h4C;
                    16'h212C: data_out = 8'h4D;
                    16'h212D: data_out = 8'h4E;
                    16'h212E: data_out = 8'h4F;
                    16'h212F: data_out = 8'h50;
                    16'h2130: data_out = 8'h51;
                    16'h2131: data_out = 8'h52;
                    16'h2132: data_out = 8'h53;
                    16'h2133: data_out = 8'h54;
                    16'h2134: data_out = 8'h55;
                    16'h2135: data_out = 8'h56;
                    16'h2136: data_out = 8'h57;
                    16'h2137: data_out = 8'h58;
                    16'h2138: data_out = 8'h59;
                    16'h2139: data_out = 8'h5A;
                    16'h213A: data_out = 8'h5B;
                    16'h213B: data_out = 8'h5C;
                    16'h213C: data_out = 8'h5D;
                    16'h213D: data_out = 8'h5E;
                    16'h213E: data_out = 8'h5F;
                    16'h213F: data_out = 8'h60;
                    16'h2140: data_out = 8'h61;
                    16'h2141: data_out = 8'h62;
                    16'h2142: data_out = 8'h63;
                    16'h2143: data_out = 8'h64;
                    16'h2144: data_out = 8'h65;
                    16'h2145: data_out = 8'h66;
                    16'h2146: data_out = 8'h67;
                    16'h2147: data_out = 8'h68;
                    16'h2148: data_out = 8'h69;
                    16'h2149: data_out = 8'h6A;
                    16'h214A: data_out = 8'h6B;
                    16'h214B: data_out = 8'h6C;
                    16'h214C: data_out = 8'h6D;
                    16'h214D: data_out = 8'h6E;
                    16'h214E: data_out = 8'h6F;
                    16'h214F: data_out = 8'h70;
                    16'h2150: data_out = 8'h71;
                    16'h2151: data_out = 8'h72;
                    16'h2152: data_out = 8'h73;
                    16'h2153: data_out = 8'h74;
                    16'h2154: data_out = 8'h75;
                    16'h2155: data_out = 8'h76;
                    16'h2156: data_out = 8'h77;
                    16'h2157: data_out = 8'h78;
                    16'h2158: data_out = 8'h79;
                    16'h2159: data_out = 8'h7A;
                    16'h215A: data_out = 8'h7B;
                    16'h215B: data_out = 8'h7C;
                    16'h215C: data_out = 8'h7D;
                    16'h215D: data_out = 8'h7E;
                    16'h215E: data_out = 8'h7F;
                    16'h215F: data_out = 8'h80;
                    16'h2160: data_out = 8'h81;
                    16'h2161: data_out = 8'h82;
                    16'h2162: data_out = 8'h83;
                    16'h2163: data_out = 8'h84;
                    16'h2164: data_out = 8'h85;
                    16'h2165: data_out = 8'h86;
                    16'h2166: data_out = 8'h87;
                    16'h2167: data_out = 8'h88;
                    16'h2168: data_out = 8'h89;
                    16'h2169: data_out = 8'h8A;
                    16'h216A: data_out = 8'h8B;
                    16'h216B: data_out = 8'h8C;
                    16'h216C: data_out = 8'h8D;
                    16'h216D: data_out = 8'h8E;
                    16'h216E: data_out = 8'h8F;
                    16'h216F: data_out = 8'h90;
                    16'h2170: data_out = 8'h91;
                    16'h2171: data_out = 8'h92;
                    16'h2172: data_out = 8'h93;
                    16'h2173: data_out = 8'h94;
                    16'h2174: data_out = 8'h95;
                    16'h2175: data_out = 8'h96;
                    16'h2176: data_out = 8'h97;
                    16'h2177: data_out = 8'h98;
                    16'h2178: data_out = 8'h99;
                    16'h2179: data_out = 8'h9A;
                    16'h217A: data_out = 8'h9B;
                    16'h217B: data_out = 8'h9C;
                    16'h217C: data_out = 8'h9D;
                    16'h217D: data_out = 8'h9E;
                    16'h217E: data_out = 8'h9F;
                    16'h217F: data_out = 8'hA0;
                    16'h2180: data_out = 8'h21;
                    16'h2181: data_out = 8'h20;
                    16'h2182: data_out = 8'h1F;
                    16'h2183: data_out = 8'h1E;
                    16'h2184: data_out = 8'h1D;
                    16'h2185: data_out = 8'h1C;
                    16'h2186: data_out = 8'h1B;
                    16'h2187: data_out = 8'h1A;
                    16'h2188: data_out = 8'h19;
                    16'h2189: data_out = 8'h18;
                    16'h218A: data_out = 8'h17;
                    16'h218B: data_out = 8'h16;
                    16'h218C: data_out = 8'h15;
                    16'h218D: data_out = 8'h14;
                    16'h218E: data_out = 8'h13;
                    16'h218F: data_out = 8'h12;
                    16'h2190: data_out = 8'h11;
                    16'h2191: data_out = 8'h10;
                    16'h2192: data_out = 8'hF;
                    16'h2193: data_out = 8'hE;
                    16'h2194: data_out = 8'hD;
                    16'h2195: data_out = 8'hC;
                    16'h2196: data_out = 8'hB;
                    16'h2197: data_out = 8'hA;
                    16'h2198: data_out = 8'h9;
                    16'h2199: data_out = 8'h8;
                    16'h219A: data_out = 8'h7;
                    16'h219B: data_out = 8'h6;
                    16'h219C: data_out = 8'h5;
                    16'h219D: data_out = 8'h4;
                    16'h219E: data_out = 8'h3;
                    16'h219F: data_out = 8'h2;
                    16'h21A0: data_out = 8'h1;
                    16'h21A1: data_out = 8'h0;
                    16'h21A2: data_out = 8'h81;
                    16'h21A3: data_out = 8'h82;
                    16'h21A4: data_out = 8'h83;
                    16'h21A5: data_out = 8'h84;
                    16'h21A6: data_out = 8'h85;
                    16'h21A7: data_out = 8'h86;
                    16'h21A8: data_out = 8'h87;
                    16'h21A9: data_out = 8'h88;
                    16'h21AA: data_out = 8'h89;
                    16'h21AB: data_out = 8'h8A;
                    16'h21AC: data_out = 8'h8B;
                    16'h21AD: data_out = 8'h8C;
                    16'h21AE: data_out = 8'h8D;
                    16'h21AF: data_out = 8'h8E;
                    16'h21B0: data_out = 8'h8F;
                    16'h21B1: data_out = 8'h90;
                    16'h21B2: data_out = 8'h91;
                    16'h21B3: data_out = 8'h92;
                    16'h21B4: data_out = 8'h93;
                    16'h21B5: data_out = 8'h94;
                    16'h21B6: data_out = 8'h95;
                    16'h21B7: data_out = 8'h96;
                    16'h21B8: data_out = 8'h97;
                    16'h21B9: data_out = 8'h98;
                    16'h21BA: data_out = 8'h99;
                    16'h21BB: data_out = 8'h9A;
                    16'h21BC: data_out = 8'h9B;
                    16'h21BD: data_out = 8'h9C;
                    16'h21BE: data_out = 8'h9D;
                    16'h21BF: data_out = 8'h9E;
                    16'h21C0: data_out = 8'h9F;
                    16'h21C1: data_out = 8'hA0;
                    16'h21C2: data_out = 8'hA1;
                    16'h21C3: data_out = 8'hA2;
                    16'h21C4: data_out = 8'hA3;
                    16'h21C5: data_out = 8'hA4;
                    16'h21C6: data_out = 8'hA5;
                    16'h21C7: data_out = 8'hA6;
                    16'h21C8: data_out = 8'hA7;
                    16'h21C9: data_out = 8'hA8;
                    16'h21CA: data_out = 8'hA9;
                    16'h21CB: data_out = 8'hAA;
                    16'h21CC: data_out = 8'hAB;
                    16'h21CD: data_out = 8'hAC;
                    16'h21CE: data_out = 8'hAD;
                    16'h21CF: data_out = 8'hAE;
                    16'h21D0: data_out = 8'hAF;
                    16'h21D1: data_out = 8'hB0;
                    16'h21D2: data_out = 8'hB1;
                    16'h21D3: data_out = 8'hB2;
                    16'h21D4: data_out = 8'hB3;
                    16'h21D5: data_out = 8'hB4;
                    16'h21D6: data_out = 8'hB5;
                    16'h21D7: data_out = 8'hB6;
                    16'h21D8: data_out = 8'hB7;
                    16'h21D9: data_out = 8'hB8;
                    16'h21DA: data_out = 8'hB9;
                    16'h21DB: data_out = 8'hBA;
                    16'h21DC: data_out = 8'hBB;
                    16'h21DD: data_out = 8'hBC;
                    16'h21DE: data_out = 8'hBD;
                    16'h21DF: data_out = 8'hBE;
                    16'h21E0: data_out = 8'hBF;
                    16'h21E1: data_out = 8'hC0;
                    16'h21E2: data_out = 8'hC1;
                    16'h21E3: data_out = 8'hC2;
                    16'h21E4: data_out = 8'hC3;
                    16'h21E5: data_out = 8'hC4;
                    16'h21E6: data_out = 8'hC5;
                    16'h21E7: data_out = 8'hC6;
                    16'h21E8: data_out = 8'hC7;
                    16'h21E9: data_out = 8'hC8;
                    16'h21EA: data_out = 8'hC9;
                    16'h21EB: data_out = 8'hCA;
                    16'h21EC: data_out = 8'hCB;
                    16'h21ED: data_out = 8'hCC;
                    16'h21EE: data_out = 8'hCD;
                    16'h21EF: data_out = 8'hCE;
                    16'h21F0: data_out = 8'hCF;
                    16'h21F1: data_out = 8'hD0;
                    16'h21F2: data_out = 8'hD1;
                    16'h21F3: data_out = 8'hD2;
                    16'h21F4: data_out = 8'hD3;
                    16'h21F5: data_out = 8'hD4;
                    16'h21F6: data_out = 8'hD5;
                    16'h21F7: data_out = 8'hD6;
                    16'h21F8: data_out = 8'hD7;
                    16'h21F9: data_out = 8'hD8;
                    16'h21FA: data_out = 8'hD9;
                    16'h21FB: data_out = 8'hDA;
                    16'h21FC: data_out = 8'hDB;
                    16'h21FD: data_out = 8'hDC;
                    16'h21FE: data_out = 8'hDD;
                    16'h21FF: data_out = 8'hDE;
                    16'h2200: data_out = 8'h22;
                    16'h2201: data_out = 8'h23;
                    16'h2202: data_out = 8'h24;
                    16'h2203: data_out = 8'h25;
                    16'h2204: data_out = 8'h26;
                    16'h2205: data_out = 8'h27;
                    16'h2206: data_out = 8'h28;
                    16'h2207: data_out = 8'h29;
                    16'h2208: data_out = 8'h2A;
                    16'h2209: data_out = 8'h2B;
                    16'h220A: data_out = 8'h2C;
                    16'h220B: data_out = 8'h2D;
                    16'h220C: data_out = 8'h2E;
                    16'h220D: data_out = 8'h2F;
                    16'h220E: data_out = 8'h30;
                    16'h220F: data_out = 8'h31;
                    16'h2210: data_out = 8'h32;
                    16'h2211: data_out = 8'h33;
                    16'h2212: data_out = 8'h34;
                    16'h2213: data_out = 8'h35;
                    16'h2214: data_out = 8'h36;
                    16'h2215: data_out = 8'h37;
                    16'h2216: data_out = 8'h38;
                    16'h2217: data_out = 8'h39;
                    16'h2218: data_out = 8'h3A;
                    16'h2219: data_out = 8'h3B;
                    16'h221A: data_out = 8'h3C;
                    16'h221B: data_out = 8'h3D;
                    16'h221C: data_out = 8'h3E;
                    16'h221D: data_out = 8'h3F;
                    16'h221E: data_out = 8'h40;
                    16'h221F: data_out = 8'h41;
                    16'h2220: data_out = 8'h42;
                    16'h2221: data_out = 8'h43;
                    16'h2222: data_out = 8'h44;
                    16'h2223: data_out = 8'h45;
                    16'h2224: data_out = 8'h46;
                    16'h2225: data_out = 8'h47;
                    16'h2226: data_out = 8'h48;
                    16'h2227: data_out = 8'h49;
                    16'h2228: data_out = 8'h4A;
                    16'h2229: data_out = 8'h4B;
                    16'h222A: data_out = 8'h4C;
                    16'h222B: data_out = 8'h4D;
                    16'h222C: data_out = 8'h4E;
                    16'h222D: data_out = 8'h4F;
                    16'h222E: data_out = 8'h50;
                    16'h222F: data_out = 8'h51;
                    16'h2230: data_out = 8'h52;
                    16'h2231: data_out = 8'h53;
                    16'h2232: data_out = 8'h54;
                    16'h2233: data_out = 8'h55;
                    16'h2234: data_out = 8'h56;
                    16'h2235: data_out = 8'h57;
                    16'h2236: data_out = 8'h58;
                    16'h2237: data_out = 8'h59;
                    16'h2238: data_out = 8'h5A;
                    16'h2239: data_out = 8'h5B;
                    16'h223A: data_out = 8'h5C;
                    16'h223B: data_out = 8'h5D;
                    16'h223C: data_out = 8'h5E;
                    16'h223D: data_out = 8'h5F;
                    16'h223E: data_out = 8'h60;
                    16'h223F: data_out = 8'h61;
                    16'h2240: data_out = 8'h62;
                    16'h2241: data_out = 8'h63;
                    16'h2242: data_out = 8'h64;
                    16'h2243: data_out = 8'h65;
                    16'h2244: data_out = 8'h66;
                    16'h2245: data_out = 8'h67;
                    16'h2246: data_out = 8'h68;
                    16'h2247: data_out = 8'h69;
                    16'h2248: data_out = 8'h6A;
                    16'h2249: data_out = 8'h6B;
                    16'h224A: data_out = 8'h6C;
                    16'h224B: data_out = 8'h6D;
                    16'h224C: data_out = 8'h6E;
                    16'h224D: data_out = 8'h6F;
                    16'h224E: data_out = 8'h70;
                    16'h224F: data_out = 8'h71;
                    16'h2250: data_out = 8'h72;
                    16'h2251: data_out = 8'h73;
                    16'h2252: data_out = 8'h74;
                    16'h2253: data_out = 8'h75;
                    16'h2254: data_out = 8'h76;
                    16'h2255: data_out = 8'h77;
                    16'h2256: data_out = 8'h78;
                    16'h2257: data_out = 8'h79;
                    16'h2258: data_out = 8'h7A;
                    16'h2259: data_out = 8'h7B;
                    16'h225A: data_out = 8'h7C;
                    16'h225B: data_out = 8'h7D;
                    16'h225C: data_out = 8'h7E;
                    16'h225D: data_out = 8'h7F;
                    16'h225E: data_out = 8'h80;
                    16'h225F: data_out = 8'h81;
                    16'h2260: data_out = 8'h82;
                    16'h2261: data_out = 8'h83;
                    16'h2262: data_out = 8'h84;
                    16'h2263: data_out = 8'h85;
                    16'h2264: data_out = 8'h86;
                    16'h2265: data_out = 8'h87;
                    16'h2266: data_out = 8'h88;
                    16'h2267: data_out = 8'h89;
                    16'h2268: data_out = 8'h8A;
                    16'h2269: data_out = 8'h8B;
                    16'h226A: data_out = 8'h8C;
                    16'h226B: data_out = 8'h8D;
                    16'h226C: data_out = 8'h8E;
                    16'h226D: data_out = 8'h8F;
                    16'h226E: data_out = 8'h90;
                    16'h226F: data_out = 8'h91;
                    16'h2270: data_out = 8'h92;
                    16'h2271: data_out = 8'h93;
                    16'h2272: data_out = 8'h94;
                    16'h2273: data_out = 8'h95;
                    16'h2274: data_out = 8'h96;
                    16'h2275: data_out = 8'h97;
                    16'h2276: data_out = 8'h98;
                    16'h2277: data_out = 8'h99;
                    16'h2278: data_out = 8'h9A;
                    16'h2279: data_out = 8'h9B;
                    16'h227A: data_out = 8'h9C;
                    16'h227B: data_out = 8'h9D;
                    16'h227C: data_out = 8'h9E;
                    16'h227D: data_out = 8'h9F;
                    16'h227E: data_out = 8'hA0;
                    16'h227F: data_out = 8'hA1;
                    16'h2280: data_out = 8'h22;
                    16'h2281: data_out = 8'h21;
                    16'h2282: data_out = 8'h20;
                    16'h2283: data_out = 8'h1F;
                    16'h2284: data_out = 8'h1E;
                    16'h2285: data_out = 8'h1D;
                    16'h2286: data_out = 8'h1C;
                    16'h2287: data_out = 8'h1B;
                    16'h2288: data_out = 8'h1A;
                    16'h2289: data_out = 8'h19;
                    16'h228A: data_out = 8'h18;
                    16'h228B: data_out = 8'h17;
                    16'h228C: data_out = 8'h16;
                    16'h228D: data_out = 8'h15;
                    16'h228E: data_out = 8'h14;
                    16'h228F: data_out = 8'h13;
                    16'h2290: data_out = 8'h12;
                    16'h2291: data_out = 8'h11;
                    16'h2292: data_out = 8'h10;
                    16'h2293: data_out = 8'hF;
                    16'h2294: data_out = 8'hE;
                    16'h2295: data_out = 8'hD;
                    16'h2296: data_out = 8'hC;
                    16'h2297: data_out = 8'hB;
                    16'h2298: data_out = 8'hA;
                    16'h2299: data_out = 8'h9;
                    16'h229A: data_out = 8'h8;
                    16'h229B: data_out = 8'h7;
                    16'h229C: data_out = 8'h6;
                    16'h229D: data_out = 8'h5;
                    16'h229E: data_out = 8'h4;
                    16'h229F: data_out = 8'h3;
                    16'h22A0: data_out = 8'h2;
                    16'h22A1: data_out = 8'h1;
                    16'h22A2: data_out = 8'h0;
                    16'h22A3: data_out = 8'h81;
                    16'h22A4: data_out = 8'h82;
                    16'h22A5: data_out = 8'h83;
                    16'h22A6: data_out = 8'h84;
                    16'h22A7: data_out = 8'h85;
                    16'h22A8: data_out = 8'h86;
                    16'h22A9: data_out = 8'h87;
                    16'h22AA: data_out = 8'h88;
                    16'h22AB: data_out = 8'h89;
                    16'h22AC: data_out = 8'h8A;
                    16'h22AD: data_out = 8'h8B;
                    16'h22AE: data_out = 8'h8C;
                    16'h22AF: data_out = 8'h8D;
                    16'h22B0: data_out = 8'h8E;
                    16'h22B1: data_out = 8'h8F;
                    16'h22B2: data_out = 8'h90;
                    16'h22B3: data_out = 8'h91;
                    16'h22B4: data_out = 8'h92;
                    16'h22B5: data_out = 8'h93;
                    16'h22B6: data_out = 8'h94;
                    16'h22B7: data_out = 8'h95;
                    16'h22B8: data_out = 8'h96;
                    16'h22B9: data_out = 8'h97;
                    16'h22BA: data_out = 8'h98;
                    16'h22BB: data_out = 8'h99;
                    16'h22BC: data_out = 8'h9A;
                    16'h22BD: data_out = 8'h9B;
                    16'h22BE: data_out = 8'h9C;
                    16'h22BF: data_out = 8'h9D;
                    16'h22C0: data_out = 8'h9E;
                    16'h22C1: data_out = 8'h9F;
                    16'h22C2: data_out = 8'hA0;
                    16'h22C3: data_out = 8'hA1;
                    16'h22C4: data_out = 8'hA2;
                    16'h22C5: data_out = 8'hA3;
                    16'h22C6: data_out = 8'hA4;
                    16'h22C7: data_out = 8'hA5;
                    16'h22C8: data_out = 8'hA6;
                    16'h22C9: data_out = 8'hA7;
                    16'h22CA: data_out = 8'hA8;
                    16'h22CB: data_out = 8'hA9;
                    16'h22CC: data_out = 8'hAA;
                    16'h22CD: data_out = 8'hAB;
                    16'h22CE: data_out = 8'hAC;
                    16'h22CF: data_out = 8'hAD;
                    16'h22D0: data_out = 8'hAE;
                    16'h22D1: data_out = 8'hAF;
                    16'h22D2: data_out = 8'hB0;
                    16'h22D3: data_out = 8'hB1;
                    16'h22D4: data_out = 8'hB2;
                    16'h22D5: data_out = 8'hB3;
                    16'h22D6: data_out = 8'hB4;
                    16'h22D7: data_out = 8'hB5;
                    16'h22D8: data_out = 8'hB6;
                    16'h22D9: data_out = 8'hB7;
                    16'h22DA: data_out = 8'hB8;
                    16'h22DB: data_out = 8'hB9;
                    16'h22DC: data_out = 8'hBA;
                    16'h22DD: data_out = 8'hBB;
                    16'h22DE: data_out = 8'hBC;
                    16'h22DF: data_out = 8'hBD;
                    16'h22E0: data_out = 8'hBE;
                    16'h22E1: data_out = 8'hBF;
                    16'h22E2: data_out = 8'hC0;
                    16'h22E3: data_out = 8'hC1;
                    16'h22E4: data_out = 8'hC2;
                    16'h22E5: data_out = 8'hC3;
                    16'h22E6: data_out = 8'hC4;
                    16'h22E7: data_out = 8'hC5;
                    16'h22E8: data_out = 8'hC6;
                    16'h22E9: data_out = 8'hC7;
                    16'h22EA: data_out = 8'hC8;
                    16'h22EB: data_out = 8'hC9;
                    16'h22EC: data_out = 8'hCA;
                    16'h22ED: data_out = 8'hCB;
                    16'h22EE: data_out = 8'hCC;
                    16'h22EF: data_out = 8'hCD;
                    16'h22F0: data_out = 8'hCE;
                    16'h22F1: data_out = 8'hCF;
                    16'h22F2: data_out = 8'hD0;
                    16'h22F3: data_out = 8'hD1;
                    16'h22F4: data_out = 8'hD2;
                    16'h22F5: data_out = 8'hD3;
                    16'h22F6: data_out = 8'hD4;
                    16'h22F7: data_out = 8'hD5;
                    16'h22F8: data_out = 8'hD6;
                    16'h22F9: data_out = 8'hD7;
                    16'h22FA: data_out = 8'hD8;
                    16'h22FB: data_out = 8'hD9;
                    16'h22FC: data_out = 8'hDA;
                    16'h22FD: data_out = 8'hDB;
                    16'h22FE: data_out = 8'hDC;
                    16'h22FF: data_out = 8'hDD;
                    16'h2300: data_out = 8'h23;
                    16'h2301: data_out = 8'h24;
                    16'h2302: data_out = 8'h25;
                    16'h2303: data_out = 8'h26;
                    16'h2304: data_out = 8'h27;
                    16'h2305: data_out = 8'h28;
                    16'h2306: data_out = 8'h29;
                    16'h2307: data_out = 8'h2A;
                    16'h2308: data_out = 8'h2B;
                    16'h2309: data_out = 8'h2C;
                    16'h230A: data_out = 8'h2D;
                    16'h230B: data_out = 8'h2E;
                    16'h230C: data_out = 8'h2F;
                    16'h230D: data_out = 8'h30;
                    16'h230E: data_out = 8'h31;
                    16'h230F: data_out = 8'h32;
                    16'h2310: data_out = 8'h33;
                    16'h2311: data_out = 8'h34;
                    16'h2312: data_out = 8'h35;
                    16'h2313: data_out = 8'h36;
                    16'h2314: data_out = 8'h37;
                    16'h2315: data_out = 8'h38;
                    16'h2316: data_out = 8'h39;
                    16'h2317: data_out = 8'h3A;
                    16'h2318: data_out = 8'h3B;
                    16'h2319: data_out = 8'h3C;
                    16'h231A: data_out = 8'h3D;
                    16'h231B: data_out = 8'h3E;
                    16'h231C: data_out = 8'h3F;
                    16'h231D: data_out = 8'h40;
                    16'h231E: data_out = 8'h41;
                    16'h231F: data_out = 8'h42;
                    16'h2320: data_out = 8'h43;
                    16'h2321: data_out = 8'h44;
                    16'h2322: data_out = 8'h45;
                    16'h2323: data_out = 8'h46;
                    16'h2324: data_out = 8'h47;
                    16'h2325: data_out = 8'h48;
                    16'h2326: data_out = 8'h49;
                    16'h2327: data_out = 8'h4A;
                    16'h2328: data_out = 8'h4B;
                    16'h2329: data_out = 8'h4C;
                    16'h232A: data_out = 8'h4D;
                    16'h232B: data_out = 8'h4E;
                    16'h232C: data_out = 8'h4F;
                    16'h232D: data_out = 8'h50;
                    16'h232E: data_out = 8'h51;
                    16'h232F: data_out = 8'h52;
                    16'h2330: data_out = 8'h53;
                    16'h2331: data_out = 8'h54;
                    16'h2332: data_out = 8'h55;
                    16'h2333: data_out = 8'h56;
                    16'h2334: data_out = 8'h57;
                    16'h2335: data_out = 8'h58;
                    16'h2336: data_out = 8'h59;
                    16'h2337: data_out = 8'h5A;
                    16'h2338: data_out = 8'h5B;
                    16'h2339: data_out = 8'h5C;
                    16'h233A: data_out = 8'h5D;
                    16'h233B: data_out = 8'h5E;
                    16'h233C: data_out = 8'h5F;
                    16'h233D: data_out = 8'h60;
                    16'h233E: data_out = 8'h61;
                    16'h233F: data_out = 8'h62;
                    16'h2340: data_out = 8'h63;
                    16'h2341: data_out = 8'h64;
                    16'h2342: data_out = 8'h65;
                    16'h2343: data_out = 8'h66;
                    16'h2344: data_out = 8'h67;
                    16'h2345: data_out = 8'h68;
                    16'h2346: data_out = 8'h69;
                    16'h2347: data_out = 8'h6A;
                    16'h2348: data_out = 8'h6B;
                    16'h2349: data_out = 8'h6C;
                    16'h234A: data_out = 8'h6D;
                    16'h234B: data_out = 8'h6E;
                    16'h234C: data_out = 8'h6F;
                    16'h234D: data_out = 8'h70;
                    16'h234E: data_out = 8'h71;
                    16'h234F: data_out = 8'h72;
                    16'h2350: data_out = 8'h73;
                    16'h2351: data_out = 8'h74;
                    16'h2352: data_out = 8'h75;
                    16'h2353: data_out = 8'h76;
                    16'h2354: data_out = 8'h77;
                    16'h2355: data_out = 8'h78;
                    16'h2356: data_out = 8'h79;
                    16'h2357: data_out = 8'h7A;
                    16'h2358: data_out = 8'h7B;
                    16'h2359: data_out = 8'h7C;
                    16'h235A: data_out = 8'h7D;
                    16'h235B: data_out = 8'h7E;
                    16'h235C: data_out = 8'h7F;
                    16'h235D: data_out = 8'h80;
                    16'h235E: data_out = 8'h81;
                    16'h235F: data_out = 8'h82;
                    16'h2360: data_out = 8'h83;
                    16'h2361: data_out = 8'h84;
                    16'h2362: data_out = 8'h85;
                    16'h2363: data_out = 8'h86;
                    16'h2364: data_out = 8'h87;
                    16'h2365: data_out = 8'h88;
                    16'h2366: data_out = 8'h89;
                    16'h2367: data_out = 8'h8A;
                    16'h2368: data_out = 8'h8B;
                    16'h2369: data_out = 8'h8C;
                    16'h236A: data_out = 8'h8D;
                    16'h236B: data_out = 8'h8E;
                    16'h236C: data_out = 8'h8F;
                    16'h236D: data_out = 8'h90;
                    16'h236E: data_out = 8'h91;
                    16'h236F: data_out = 8'h92;
                    16'h2370: data_out = 8'h93;
                    16'h2371: data_out = 8'h94;
                    16'h2372: data_out = 8'h95;
                    16'h2373: data_out = 8'h96;
                    16'h2374: data_out = 8'h97;
                    16'h2375: data_out = 8'h98;
                    16'h2376: data_out = 8'h99;
                    16'h2377: data_out = 8'h9A;
                    16'h2378: data_out = 8'h9B;
                    16'h2379: data_out = 8'h9C;
                    16'h237A: data_out = 8'h9D;
                    16'h237B: data_out = 8'h9E;
                    16'h237C: data_out = 8'h9F;
                    16'h237D: data_out = 8'hA0;
                    16'h237E: data_out = 8'hA1;
                    16'h237F: data_out = 8'hA2;
                    16'h2380: data_out = 8'h23;
                    16'h2381: data_out = 8'h22;
                    16'h2382: data_out = 8'h21;
                    16'h2383: data_out = 8'h20;
                    16'h2384: data_out = 8'h1F;
                    16'h2385: data_out = 8'h1E;
                    16'h2386: data_out = 8'h1D;
                    16'h2387: data_out = 8'h1C;
                    16'h2388: data_out = 8'h1B;
                    16'h2389: data_out = 8'h1A;
                    16'h238A: data_out = 8'h19;
                    16'h238B: data_out = 8'h18;
                    16'h238C: data_out = 8'h17;
                    16'h238D: data_out = 8'h16;
                    16'h238E: data_out = 8'h15;
                    16'h238F: data_out = 8'h14;
                    16'h2390: data_out = 8'h13;
                    16'h2391: data_out = 8'h12;
                    16'h2392: data_out = 8'h11;
                    16'h2393: data_out = 8'h10;
                    16'h2394: data_out = 8'hF;
                    16'h2395: data_out = 8'hE;
                    16'h2396: data_out = 8'hD;
                    16'h2397: data_out = 8'hC;
                    16'h2398: data_out = 8'hB;
                    16'h2399: data_out = 8'hA;
                    16'h239A: data_out = 8'h9;
                    16'h239B: data_out = 8'h8;
                    16'h239C: data_out = 8'h7;
                    16'h239D: data_out = 8'h6;
                    16'h239E: data_out = 8'h5;
                    16'h239F: data_out = 8'h4;
                    16'h23A0: data_out = 8'h3;
                    16'h23A1: data_out = 8'h2;
                    16'h23A2: data_out = 8'h1;
                    16'h23A3: data_out = 8'h0;
                    16'h23A4: data_out = 8'h81;
                    16'h23A5: data_out = 8'h82;
                    16'h23A6: data_out = 8'h83;
                    16'h23A7: data_out = 8'h84;
                    16'h23A8: data_out = 8'h85;
                    16'h23A9: data_out = 8'h86;
                    16'h23AA: data_out = 8'h87;
                    16'h23AB: data_out = 8'h88;
                    16'h23AC: data_out = 8'h89;
                    16'h23AD: data_out = 8'h8A;
                    16'h23AE: data_out = 8'h8B;
                    16'h23AF: data_out = 8'h8C;
                    16'h23B0: data_out = 8'h8D;
                    16'h23B1: data_out = 8'h8E;
                    16'h23B2: data_out = 8'h8F;
                    16'h23B3: data_out = 8'h90;
                    16'h23B4: data_out = 8'h91;
                    16'h23B5: data_out = 8'h92;
                    16'h23B6: data_out = 8'h93;
                    16'h23B7: data_out = 8'h94;
                    16'h23B8: data_out = 8'h95;
                    16'h23B9: data_out = 8'h96;
                    16'h23BA: data_out = 8'h97;
                    16'h23BB: data_out = 8'h98;
                    16'h23BC: data_out = 8'h99;
                    16'h23BD: data_out = 8'h9A;
                    16'h23BE: data_out = 8'h9B;
                    16'h23BF: data_out = 8'h9C;
                    16'h23C0: data_out = 8'h9D;
                    16'h23C1: data_out = 8'h9E;
                    16'h23C2: data_out = 8'h9F;
                    16'h23C3: data_out = 8'hA0;
                    16'h23C4: data_out = 8'hA1;
                    16'h23C5: data_out = 8'hA2;
                    16'h23C6: data_out = 8'hA3;
                    16'h23C7: data_out = 8'hA4;
                    16'h23C8: data_out = 8'hA5;
                    16'h23C9: data_out = 8'hA6;
                    16'h23CA: data_out = 8'hA7;
                    16'h23CB: data_out = 8'hA8;
                    16'h23CC: data_out = 8'hA9;
                    16'h23CD: data_out = 8'hAA;
                    16'h23CE: data_out = 8'hAB;
                    16'h23CF: data_out = 8'hAC;
                    16'h23D0: data_out = 8'hAD;
                    16'h23D1: data_out = 8'hAE;
                    16'h23D2: data_out = 8'hAF;
                    16'h23D3: data_out = 8'hB0;
                    16'h23D4: data_out = 8'hB1;
                    16'h23D5: data_out = 8'hB2;
                    16'h23D6: data_out = 8'hB3;
                    16'h23D7: data_out = 8'hB4;
                    16'h23D8: data_out = 8'hB5;
                    16'h23D9: data_out = 8'hB6;
                    16'h23DA: data_out = 8'hB7;
                    16'h23DB: data_out = 8'hB8;
                    16'h23DC: data_out = 8'hB9;
                    16'h23DD: data_out = 8'hBA;
                    16'h23DE: data_out = 8'hBB;
                    16'h23DF: data_out = 8'hBC;
                    16'h23E0: data_out = 8'hBD;
                    16'h23E1: data_out = 8'hBE;
                    16'h23E2: data_out = 8'hBF;
                    16'h23E3: data_out = 8'hC0;
                    16'h23E4: data_out = 8'hC1;
                    16'h23E5: data_out = 8'hC2;
                    16'h23E6: data_out = 8'hC3;
                    16'h23E7: data_out = 8'hC4;
                    16'h23E8: data_out = 8'hC5;
                    16'h23E9: data_out = 8'hC6;
                    16'h23EA: data_out = 8'hC7;
                    16'h23EB: data_out = 8'hC8;
                    16'h23EC: data_out = 8'hC9;
                    16'h23ED: data_out = 8'hCA;
                    16'h23EE: data_out = 8'hCB;
                    16'h23EF: data_out = 8'hCC;
                    16'h23F0: data_out = 8'hCD;
                    16'h23F1: data_out = 8'hCE;
                    16'h23F2: data_out = 8'hCF;
                    16'h23F3: data_out = 8'hD0;
                    16'h23F4: data_out = 8'hD1;
                    16'h23F5: data_out = 8'hD2;
                    16'h23F6: data_out = 8'hD3;
                    16'h23F7: data_out = 8'hD4;
                    16'h23F8: data_out = 8'hD5;
                    16'h23F9: data_out = 8'hD6;
                    16'h23FA: data_out = 8'hD7;
                    16'h23FB: data_out = 8'hD8;
                    16'h23FC: data_out = 8'hD9;
                    16'h23FD: data_out = 8'hDA;
                    16'h23FE: data_out = 8'hDB;
                    16'h23FF: data_out = 8'hDC;
                    16'h2400: data_out = 8'h24;
                    16'h2401: data_out = 8'h25;
                    16'h2402: data_out = 8'h26;
                    16'h2403: data_out = 8'h27;
                    16'h2404: data_out = 8'h28;
                    16'h2405: data_out = 8'h29;
                    16'h2406: data_out = 8'h2A;
                    16'h2407: data_out = 8'h2B;
                    16'h2408: data_out = 8'h2C;
                    16'h2409: data_out = 8'h2D;
                    16'h240A: data_out = 8'h2E;
                    16'h240B: data_out = 8'h2F;
                    16'h240C: data_out = 8'h30;
                    16'h240D: data_out = 8'h31;
                    16'h240E: data_out = 8'h32;
                    16'h240F: data_out = 8'h33;
                    16'h2410: data_out = 8'h34;
                    16'h2411: data_out = 8'h35;
                    16'h2412: data_out = 8'h36;
                    16'h2413: data_out = 8'h37;
                    16'h2414: data_out = 8'h38;
                    16'h2415: data_out = 8'h39;
                    16'h2416: data_out = 8'h3A;
                    16'h2417: data_out = 8'h3B;
                    16'h2418: data_out = 8'h3C;
                    16'h2419: data_out = 8'h3D;
                    16'h241A: data_out = 8'h3E;
                    16'h241B: data_out = 8'h3F;
                    16'h241C: data_out = 8'h40;
                    16'h241D: data_out = 8'h41;
                    16'h241E: data_out = 8'h42;
                    16'h241F: data_out = 8'h43;
                    16'h2420: data_out = 8'h44;
                    16'h2421: data_out = 8'h45;
                    16'h2422: data_out = 8'h46;
                    16'h2423: data_out = 8'h47;
                    16'h2424: data_out = 8'h48;
                    16'h2425: data_out = 8'h49;
                    16'h2426: data_out = 8'h4A;
                    16'h2427: data_out = 8'h4B;
                    16'h2428: data_out = 8'h4C;
                    16'h2429: data_out = 8'h4D;
                    16'h242A: data_out = 8'h4E;
                    16'h242B: data_out = 8'h4F;
                    16'h242C: data_out = 8'h50;
                    16'h242D: data_out = 8'h51;
                    16'h242E: data_out = 8'h52;
                    16'h242F: data_out = 8'h53;
                    16'h2430: data_out = 8'h54;
                    16'h2431: data_out = 8'h55;
                    16'h2432: data_out = 8'h56;
                    16'h2433: data_out = 8'h57;
                    16'h2434: data_out = 8'h58;
                    16'h2435: data_out = 8'h59;
                    16'h2436: data_out = 8'h5A;
                    16'h2437: data_out = 8'h5B;
                    16'h2438: data_out = 8'h5C;
                    16'h2439: data_out = 8'h5D;
                    16'h243A: data_out = 8'h5E;
                    16'h243B: data_out = 8'h5F;
                    16'h243C: data_out = 8'h60;
                    16'h243D: data_out = 8'h61;
                    16'h243E: data_out = 8'h62;
                    16'h243F: data_out = 8'h63;
                    16'h2440: data_out = 8'h64;
                    16'h2441: data_out = 8'h65;
                    16'h2442: data_out = 8'h66;
                    16'h2443: data_out = 8'h67;
                    16'h2444: data_out = 8'h68;
                    16'h2445: data_out = 8'h69;
                    16'h2446: data_out = 8'h6A;
                    16'h2447: data_out = 8'h6B;
                    16'h2448: data_out = 8'h6C;
                    16'h2449: data_out = 8'h6D;
                    16'h244A: data_out = 8'h6E;
                    16'h244B: data_out = 8'h6F;
                    16'h244C: data_out = 8'h70;
                    16'h244D: data_out = 8'h71;
                    16'h244E: data_out = 8'h72;
                    16'h244F: data_out = 8'h73;
                    16'h2450: data_out = 8'h74;
                    16'h2451: data_out = 8'h75;
                    16'h2452: data_out = 8'h76;
                    16'h2453: data_out = 8'h77;
                    16'h2454: data_out = 8'h78;
                    16'h2455: data_out = 8'h79;
                    16'h2456: data_out = 8'h7A;
                    16'h2457: data_out = 8'h7B;
                    16'h2458: data_out = 8'h7C;
                    16'h2459: data_out = 8'h7D;
                    16'h245A: data_out = 8'h7E;
                    16'h245B: data_out = 8'h7F;
                    16'h245C: data_out = 8'h80;
                    16'h245D: data_out = 8'h81;
                    16'h245E: data_out = 8'h82;
                    16'h245F: data_out = 8'h83;
                    16'h2460: data_out = 8'h84;
                    16'h2461: data_out = 8'h85;
                    16'h2462: data_out = 8'h86;
                    16'h2463: data_out = 8'h87;
                    16'h2464: data_out = 8'h88;
                    16'h2465: data_out = 8'h89;
                    16'h2466: data_out = 8'h8A;
                    16'h2467: data_out = 8'h8B;
                    16'h2468: data_out = 8'h8C;
                    16'h2469: data_out = 8'h8D;
                    16'h246A: data_out = 8'h8E;
                    16'h246B: data_out = 8'h8F;
                    16'h246C: data_out = 8'h90;
                    16'h246D: data_out = 8'h91;
                    16'h246E: data_out = 8'h92;
                    16'h246F: data_out = 8'h93;
                    16'h2470: data_out = 8'h94;
                    16'h2471: data_out = 8'h95;
                    16'h2472: data_out = 8'h96;
                    16'h2473: data_out = 8'h97;
                    16'h2474: data_out = 8'h98;
                    16'h2475: data_out = 8'h99;
                    16'h2476: data_out = 8'h9A;
                    16'h2477: data_out = 8'h9B;
                    16'h2478: data_out = 8'h9C;
                    16'h2479: data_out = 8'h9D;
                    16'h247A: data_out = 8'h9E;
                    16'h247B: data_out = 8'h9F;
                    16'h247C: data_out = 8'hA0;
                    16'h247D: data_out = 8'hA1;
                    16'h247E: data_out = 8'hA2;
                    16'h247F: data_out = 8'hA3;
                    16'h2480: data_out = 8'h24;
                    16'h2481: data_out = 8'h23;
                    16'h2482: data_out = 8'h22;
                    16'h2483: data_out = 8'h21;
                    16'h2484: data_out = 8'h20;
                    16'h2485: data_out = 8'h1F;
                    16'h2486: data_out = 8'h1E;
                    16'h2487: data_out = 8'h1D;
                    16'h2488: data_out = 8'h1C;
                    16'h2489: data_out = 8'h1B;
                    16'h248A: data_out = 8'h1A;
                    16'h248B: data_out = 8'h19;
                    16'h248C: data_out = 8'h18;
                    16'h248D: data_out = 8'h17;
                    16'h248E: data_out = 8'h16;
                    16'h248F: data_out = 8'h15;
                    16'h2490: data_out = 8'h14;
                    16'h2491: data_out = 8'h13;
                    16'h2492: data_out = 8'h12;
                    16'h2493: data_out = 8'h11;
                    16'h2494: data_out = 8'h10;
                    16'h2495: data_out = 8'hF;
                    16'h2496: data_out = 8'hE;
                    16'h2497: data_out = 8'hD;
                    16'h2498: data_out = 8'hC;
                    16'h2499: data_out = 8'hB;
                    16'h249A: data_out = 8'hA;
                    16'h249B: data_out = 8'h9;
                    16'h249C: data_out = 8'h8;
                    16'h249D: data_out = 8'h7;
                    16'h249E: data_out = 8'h6;
                    16'h249F: data_out = 8'h5;
                    16'h24A0: data_out = 8'h4;
                    16'h24A1: data_out = 8'h3;
                    16'h24A2: data_out = 8'h2;
                    16'h24A3: data_out = 8'h1;
                    16'h24A4: data_out = 8'h0;
                    16'h24A5: data_out = 8'h81;
                    16'h24A6: data_out = 8'h82;
                    16'h24A7: data_out = 8'h83;
                    16'h24A8: data_out = 8'h84;
                    16'h24A9: data_out = 8'h85;
                    16'h24AA: data_out = 8'h86;
                    16'h24AB: data_out = 8'h87;
                    16'h24AC: data_out = 8'h88;
                    16'h24AD: data_out = 8'h89;
                    16'h24AE: data_out = 8'h8A;
                    16'h24AF: data_out = 8'h8B;
                    16'h24B0: data_out = 8'h8C;
                    16'h24B1: data_out = 8'h8D;
                    16'h24B2: data_out = 8'h8E;
                    16'h24B3: data_out = 8'h8F;
                    16'h24B4: data_out = 8'h90;
                    16'h24B5: data_out = 8'h91;
                    16'h24B6: data_out = 8'h92;
                    16'h24B7: data_out = 8'h93;
                    16'h24B8: data_out = 8'h94;
                    16'h24B9: data_out = 8'h95;
                    16'h24BA: data_out = 8'h96;
                    16'h24BB: data_out = 8'h97;
                    16'h24BC: data_out = 8'h98;
                    16'h24BD: data_out = 8'h99;
                    16'h24BE: data_out = 8'h9A;
                    16'h24BF: data_out = 8'h9B;
                    16'h24C0: data_out = 8'h9C;
                    16'h24C1: data_out = 8'h9D;
                    16'h24C2: data_out = 8'h9E;
                    16'h24C3: data_out = 8'h9F;
                    16'h24C4: data_out = 8'hA0;
                    16'h24C5: data_out = 8'hA1;
                    16'h24C6: data_out = 8'hA2;
                    16'h24C7: data_out = 8'hA3;
                    16'h24C8: data_out = 8'hA4;
                    16'h24C9: data_out = 8'hA5;
                    16'h24CA: data_out = 8'hA6;
                    16'h24CB: data_out = 8'hA7;
                    16'h24CC: data_out = 8'hA8;
                    16'h24CD: data_out = 8'hA9;
                    16'h24CE: data_out = 8'hAA;
                    16'h24CF: data_out = 8'hAB;
                    16'h24D0: data_out = 8'hAC;
                    16'h24D1: data_out = 8'hAD;
                    16'h24D2: data_out = 8'hAE;
                    16'h24D3: data_out = 8'hAF;
                    16'h24D4: data_out = 8'hB0;
                    16'h24D5: data_out = 8'hB1;
                    16'h24D6: data_out = 8'hB2;
                    16'h24D7: data_out = 8'hB3;
                    16'h24D8: data_out = 8'hB4;
                    16'h24D9: data_out = 8'hB5;
                    16'h24DA: data_out = 8'hB6;
                    16'h24DB: data_out = 8'hB7;
                    16'h24DC: data_out = 8'hB8;
                    16'h24DD: data_out = 8'hB9;
                    16'h24DE: data_out = 8'hBA;
                    16'h24DF: data_out = 8'hBB;
                    16'h24E0: data_out = 8'hBC;
                    16'h24E1: data_out = 8'hBD;
                    16'h24E2: data_out = 8'hBE;
                    16'h24E3: data_out = 8'hBF;
                    16'h24E4: data_out = 8'hC0;
                    16'h24E5: data_out = 8'hC1;
                    16'h24E6: data_out = 8'hC2;
                    16'h24E7: data_out = 8'hC3;
                    16'h24E8: data_out = 8'hC4;
                    16'h24E9: data_out = 8'hC5;
                    16'h24EA: data_out = 8'hC6;
                    16'h24EB: data_out = 8'hC7;
                    16'h24EC: data_out = 8'hC8;
                    16'h24ED: data_out = 8'hC9;
                    16'h24EE: data_out = 8'hCA;
                    16'h24EF: data_out = 8'hCB;
                    16'h24F0: data_out = 8'hCC;
                    16'h24F1: data_out = 8'hCD;
                    16'h24F2: data_out = 8'hCE;
                    16'h24F3: data_out = 8'hCF;
                    16'h24F4: data_out = 8'hD0;
                    16'h24F5: data_out = 8'hD1;
                    16'h24F6: data_out = 8'hD2;
                    16'h24F7: data_out = 8'hD3;
                    16'h24F8: data_out = 8'hD4;
                    16'h24F9: data_out = 8'hD5;
                    16'h24FA: data_out = 8'hD6;
                    16'h24FB: data_out = 8'hD7;
                    16'h24FC: data_out = 8'hD8;
                    16'h24FD: data_out = 8'hD9;
                    16'h24FE: data_out = 8'hDA;
                    16'h24FF: data_out = 8'hDB;
                    16'h2500: data_out = 8'h25;
                    16'h2501: data_out = 8'h26;
                    16'h2502: data_out = 8'h27;
                    16'h2503: data_out = 8'h28;
                    16'h2504: data_out = 8'h29;
                    16'h2505: data_out = 8'h2A;
                    16'h2506: data_out = 8'h2B;
                    16'h2507: data_out = 8'h2C;
                    16'h2508: data_out = 8'h2D;
                    16'h2509: data_out = 8'h2E;
                    16'h250A: data_out = 8'h2F;
                    16'h250B: data_out = 8'h30;
                    16'h250C: data_out = 8'h31;
                    16'h250D: data_out = 8'h32;
                    16'h250E: data_out = 8'h33;
                    16'h250F: data_out = 8'h34;
                    16'h2510: data_out = 8'h35;
                    16'h2511: data_out = 8'h36;
                    16'h2512: data_out = 8'h37;
                    16'h2513: data_out = 8'h38;
                    16'h2514: data_out = 8'h39;
                    16'h2515: data_out = 8'h3A;
                    16'h2516: data_out = 8'h3B;
                    16'h2517: data_out = 8'h3C;
                    16'h2518: data_out = 8'h3D;
                    16'h2519: data_out = 8'h3E;
                    16'h251A: data_out = 8'h3F;
                    16'h251B: data_out = 8'h40;
                    16'h251C: data_out = 8'h41;
                    16'h251D: data_out = 8'h42;
                    16'h251E: data_out = 8'h43;
                    16'h251F: data_out = 8'h44;
                    16'h2520: data_out = 8'h45;
                    16'h2521: data_out = 8'h46;
                    16'h2522: data_out = 8'h47;
                    16'h2523: data_out = 8'h48;
                    16'h2524: data_out = 8'h49;
                    16'h2525: data_out = 8'h4A;
                    16'h2526: data_out = 8'h4B;
                    16'h2527: data_out = 8'h4C;
                    16'h2528: data_out = 8'h4D;
                    16'h2529: data_out = 8'h4E;
                    16'h252A: data_out = 8'h4F;
                    16'h252B: data_out = 8'h50;
                    16'h252C: data_out = 8'h51;
                    16'h252D: data_out = 8'h52;
                    16'h252E: data_out = 8'h53;
                    16'h252F: data_out = 8'h54;
                    16'h2530: data_out = 8'h55;
                    16'h2531: data_out = 8'h56;
                    16'h2532: data_out = 8'h57;
                    16'h2533: data_out = 8'h58;
                    16'h2534: data_out = 8'h59;
                    16'h2535: data_out = 8'h5A;
                    16'h2536: data_out = 8'h5B;
                    16'h2537: data_out = 8'h5C;
                    16'h2538: data_out = 8'h5D;
                    16'h2539: data_out = 8'h5E;
                    16'h253A: data_out = 8'h5F;
                    16'h253B: data_out = 8'h60;
                    16'h253C: data_out = 8'h61;
                    16'h253D: data_out = 8'h62;
                    16'h253E: data_out = 8'h63;
                    16'h253F: data_out = 8'h64;
                    16'h2540: data_out = 8'h65;
                    16'h2541: data_out = 8'h66;
                    16'h2542: data_out = 8'h67;
                    16'h2543: data_out = 8'h68;
                    16'h2544: data_out = 8'h69;
                    16'h2545: data_out = 8'h6A;
                    16'h2546: data_out = 8'h6B;
                    16'h2547: data_out = 8'h6C;
                    16'h2548: data_out = 8'h6D;
                    16'h2549: data_out = 8'h6E;
                    16'h254A: data_out = 8'h6F;
                    16'h254B: data_out = 8'h70;
                    16'h254C: data_out = 8'h71;
                    16'h254D: data_out = 8'h72;
                    16'h254E: data_out = 8'h73;
                    16'h254F: data_out = 8'h74;
                    16'h2550: data_out = 8'h75;
                    16'h2551: data_out = 8'h76;
                    16'h2552: data_out = 8'h77;
                    16'h2553: data_out = 8'h78;
                    16'h2554: data_out = 8'h79;
                    16'h2555: data_out = 8'h7A;
                    16'h2556: data_out = 8'h7B;
                    16'h2557: data_out = 8'h7C;
                    16'h2558: data_out = 8'h7D;
                    16'h2559: data_out = 8'h7E;
                    16'h255A: data_out = 8'h7F;
                    16'h255B: data_out = 8'h80;
                    16'h255C: data_out = 8'h81;
                    16'h255D: data_out = 8'h82;
                    16'h255E: data_out = 8'h83;
                    16'h255F: data_out = 8'h84;
                    16'h2560: data_out = 8'h85;
                    16'h2561: data_out = 8'h86;
                    16'h2562: data_out = 8'h87;
                    16'h2563: data_out = 8'h88;
                    16'h2564: data_out = 8'h89;
                    16'h2565: data_out = 8'h8A;
                    16'h2566: data_out = 8'h8B;
                    16'h2567: data_out = 8'h8C;
                    16'h2568: data_out = 8'h8D;
                    16'h2569: data_out = 8'h8E;
                    16'h256A: data_out = 8'h8F;
                    16'h256B: data_out = 8'h90;
                    16'h256C: data_out = 8'h91;
                    16'h256D: data_out = 8'h92;
                    16'h256E: data_out = 8'h93;
                    16'h256F: data_out = 8'h94;
                    16'h2570: data_out = 8'h95;
                    16'h2571: data_out = 8'h96;
                    16'h2572: data_out = 8'h97;
                    16'h2573: data_out = 8'h98;
                    16'h2574: data_out = 8'h99;
                    16'h2575: data_out = 8'h9A;
                    16'h2576: data_out = 8'h9B;
                    16'h2577: data_out = 8'h9C;
                    16'h2578: data_out = 8'h9D;
                    16'h2579: data_out = 8'h9E;
                    16'h257A: data_out = 8'h9F;
                    16'h257B: data_out = 8'hA0;
                    16'h257C: data_out = 8'hA1;
                    16'h257D: data_out = 8'hA2;
                    16'h257E: data_out = 8'hA3;
                    16'h257F: data_out = 8'hA4;
                    16'h2580: data_out = 8'h25;
                    16'h2581: data_out = 8'h24;
                    16'h2582: data_out = 8'h23;
                    16'h2583: data_out = 8'h22;
                    16'h2584: data_out = 8'h21;
                    16'h2585: data_out = 8'h20;
                    16'h2586: data_out = 8'h1F;
                    16'h2587: data_out = 8'h1E;
                    16'h2588: data_out = 8'h1D;
                    16'h2589: data_out = 8'h1C;
                    16'h258A: data_out = 8'h1B;
                    16'h258B: data_out = 8'h1A;
                    16'h258C: data_out = 8'h19;
                    16'h258D: data_out = 8'h18;
                    16'h258E: data_out = 8'h17;
                    16'h258F: data_out = 8'h16;
                    16'h2590: data_out = 8'h15;
                    16'h2591: data_out = 8'h14;
                    16'h2592: data_out = 8'h13;
                    16'h2593: data_out = 8'h12;
                    16'h2594: data_out = 8'h11;
                    16'h2595: data_out = 8'h10;
                    16'h2596: data_out = 8'hF;
                    16'h2597: data_out = 8'hE;
                    16'h2598: data_out = 8'hD;
                    16'h2599: data_out = 8'hC;
                    16'h259A: data_out = 8'hB;
                    16'h259B: data_out = 8'hA;
                    16'h259C: data_out = 8'h9;
                    16'h259D: data_out = 8'h8;
                    16'h259E: data_out = 8'h7;
                    16'h259F: data_out = 8'h6;
                    16'h25A0: data_out = 8'h5;
                    16'h25A1: data_out = 8'h4;
                    16'h25A2: data_out = 8'h3;
                    16'h25A3: data_out = 8'h2;
                    16'h25A4: data_out = 8'h1;
                    16'h25A5: data_out = 8'h0;
                    16'h25A6: data_out = 8'h81;
                    16'h25A7: data_out = 8'h82;
                    16'h25A8: data_out = 8'h83;
                    16'h25A9: data_out = 8'h84;
                    16'h25AA: data_out = 8'h85;
                    16'h25AB: data_out = 8'h86;
                    16'h25AC: data_out = 8'h87;
                    16'h25AD: data_out = 8'h88;
                    16'h25AE: data_out = 8'h89;
                    16'h25AF: data_out = 8'h8A;
                    16'h25B0: data_out = 8'h8B;
                    16'h25B1: data_out = 8'h8C;
                    16'h25B2: data_out = 8'h8D;
                    16'h25B3: data_out = 8'h8E;
                    16'h25B4: data_out = 8'h8F;
                    16'h25B5: data_out = 8'h90;
                    16'h25B6: data_out = 8'h91;
                    16'h25B7: data_out = 8'h92;
                    16'h25B8: data_out = 8'h93;
                    16'h25B9: data_out = 8'h94;
                    16'h25BA: data_out = 8'h95;
                    16'h25BB: data_out = 8'h96;
                    16'h25BC: data_out = 8'h97;
                    16'h25BD: data_out = 8'h98;
                    16'h25BE: data_out = 8'h99;
                    16'h25BF: data_out = 8'h9A;
                    16'h25C0: data_out = 8'h9B;
                    16'h25C1: data_out = 8'h9C;
                    16'h25C2: data_out = 8'h9D;
                    16'h25C3: data_out = 8'h9E;
                    16'h25C4: data_out = 8'h9F;
                    16'h25C5: data_out = 8'hA0;
                    16'h25C6: data_out = 8'hA1;
                    16'h25C7: data_out = 8'hA2;
                    16'h25C8: data_out = 8'hA3;
                    16'h25C9: data_out = 8'hA4;
                    16'h25CA: data_out = 8'hA5;
                    16'h25CB: data_out = 8'hA6;
                    16'h25CC: data_out = 8'hA7;
                    16'h25CD: data_out = 8'hA8;
                    16'h25CE: data_out = 8'hA9;
                    16'h25CF: data_out = 8'hAA;
                    16'h25D0: data_out = 8'hAB;
                    16'h25D1: data_out = 8'hAC;
                    16'h25D2: data_out = 8'hAD;
                    16'h25D3: data_out = 8'hAE;
                    16'h25D4: data_out = 8'hAF;
                    16'h25D5: data_out = 8'hB0;
                    16'h25D6: data_out = 8'hB1;
                    16'h25D7: data_out = 8'hB2;
                    16'h25D8: data_out = 8'hB3;
                    16'h25D9: data_out = 8'hB4;
                    16'h25DA: data_out = 8'hB5;
                    16'h25DB: data_out = 8'hB6;
                    16'h25DC: data_out = 8'hB7;
                    16'h25DD: data_out = 8'hB8;
                    16'h25DE: data_out = 8'hB9;
                    16'h25DF: data_out = 8'hBA;
                    16'h25E0: data_out = 8'hBB;
                    16'h25E1: data_out = 8'hBC;
                    16'h25E2: data_out = 8'hBD;
                    16'h25E3: data_out = 8'hBE;
                    16'h25E4: data_out = 8'hBF;
                    16'h25E5: data_out = 8'hC0;
                    16'h25E6: data_out = 8'hC1;
                    16'h25E7: data_out = 8'hC2;
                    16'h25E8: data_out = 8'hC3;
                    16'h25E9: data_out = 8'hC4;
                    16'h25EA: data_out = 8'hC5;
                    16'h25EB: data_out = 8'hC6;
                    16'h25EC: data_out = 8'hC7;
                    16'h25ED: data_out = 8'hC8;
                    16'h25EE: data_out = 8'hC9;
                    16'h25EF: data_out = 8'hCA;
                    16'h25F0: data_out = 8'hCB;
                    16'h25F1: data_out = 8'hCC;
                    16'h25F2: data_out = 8'hCD;
                    16'h25F3: data_out = 8'hCE;
                    16'h25F4: data_out = 8'hCF;
                    16'h25F5: data_out = 8'hD0;
                    16'h25F6: data_out = 8'hD1;
                    16'h25F7: data_out = 8'hD2;
                    16'h25F8: data_out = 8'hD3;
                    16'h25F9: data_out = 8'hD4;
                    16'h25FA: data_out = 8'hD5;
                    16'h25FB: data_out = 8'hD6;
                    16'h25FC: data_out = 8'hD7;
                    16'h25FD: data_out = 8'hD8;
                    16'h25FE: data_out = 8'hD9;
                    16'h25FF: data_out = 8'hDA;
                    16'h2600: data_out = 8'h26;
                    16'h2601: data_out = 8'h27;
                    16'h2602: data_out = 8'h28;
                    16'h2603: data_out = 8'h29;
                    16'h2604: data_out = 8'h2A;
                    16'h2605: data_out = 8'h2B;
                    16'h2606: data_out = 8'h2C;
                    16'h2607: data_out = 8'h2D;
                    16'h2608: data_out = 8'h2E;
                    16'h2609: data_out = 8'h2F;
                    16'h260A: data_out = 8'h30;
                    16'h260B: data_out = 8'h31;
                    16'h260C: data_out = 8'h32;
                    16'h260D: data_out = 8'h33;
                    16'h260E: data_out = 8'h34;
                    16'h260F: data_out = 8'h35;
                    16'h2610: data_out = 8'h36;
                    16'h2611: data_out = 8'h37;
                    16'h2612: data_out = 8'h38;
                    16'h2613: data_out = 8'h39;
                    16'h2614: data_out = 8'h3A;
                    16'h2615: data_out = 8'h3B;
                    16'h2616: data_out = 8'h3C;
                    16'h2617: data_out = 8'h3D;
                    16'h2618: data_out = 8'h3E;
                    16'h2619: data_out = 8'h3F;
                    16'h261A: data_out = 8'h40;
                    16'h261B: data_out = 8'h41;
                    16'h261C: data_out = 8'h42;
                    16'h261D: data_out = 8'h43;
                    16'h261E: data_out = 8'h44;
                    16'h261F: data_out = 8'h45;
                    16'h2620: data_out = 8'h46;
                    16'h2621: data_out = 8'h47;
                    16'h2622: data_out = 8'h48;
                    16'h2623: data_out = 8'h49;
                    16'h2624: data_out = 8'h4A;
                    16'h2625: data_out = 8'h4B;
                    16'h2626: data_out = 8'h4C;
                    16'h2627: data_out = 8'h4D;
                    16'h2628: data_out = 8'h4E;
                    16'h2629: data_out = 8'h4F;
                    16'h262A: data_out = 8'h50;
                    16'h262B: data_out = 8'h51;
                    16'h262C: data_out = 8'h52;
                    16'h262D: data_out = 8'h53;
                    16'h262E: data_out = 8'h54;
                    16'h262F: data_out = 8'h55;
                    16'h2630: data_out = 8'h56;
                    16'h2631: data_out = 8'h57;
                    16'h2632: data_out = 8'h58;
                    16'h2633: data_out = 8'h59;
                    16'h2634: data_out = 8'h5A;
                    16'h2635: data_out = 8'h5B;
                    16'h2636: data_out = 8'h5C;
                    16'h2637: data_out = 8'h5D;
                    16'h2638: data_out = 8'h5E;
                    16'h2639: data_out = 8'h5F;
                    16'h263A: data_out = 8'h60;
                    16'h263B: data_out = 8'h61;
                    16'h263C: data_out = 8'h62;
                    16'h263D: data_out = 8'h63;
                    16'h263E: data_out = 8'h64;
                    16'h263F: data_out = 8'h65;
                    16'h2640: data_out = 8'h66;
                    16'h2641: data_out = 8'h67;
                    16'h2642: data_out = 8'h68;
                    16'h2643: data_out = 8'h69;
                    16'h2644: data_out = 8'h6A;
                    16'h2645: data_out = 8'h6B;
                    16'h2646: data_out = 8'h6C;
                    16'h2647: data_out = 8'h6D;
                    16'h2648: data_out = 8'h6E;
                    16'h2649: data_out = 8'h6F;
                    16'h264A: data_out = 8'h70;
                    16'h264B: data_out = 8'h71;
                    16'h264C: data_out = 8'h72;
                    16'h264D: data_out = 8'h73;
                    16'h264E: data_out = 8'h74;
                    16'h264F: data_out = 8'h75;
                    16'h2650: data_out = 8'h76;
                    16'h2651: data_out = 8'h77;
                    16'h2652: data_out = 8'h78;
                    16'h2653: data_out = 8'h79;
                    16'h2654: data_out = 8'h7A;
                    16'h2655: data_out = 8'h7B;
                    16'h2656: data_out = 8'h7C;
                    16'h2657: data_out = 8'h7D;
                    16'h2658: data_out = 8'h7E;
                    16'h2659: data_out = 8'h7F;
                    16'h265A: data_out = 8'h80;
                    16'h265B: data_out = 8'h81;
                    16'h265C: data_out = 8'h82;
                    16'h265D: data_out = 8'h83;
                    16'h265E: data_out = 8'h84;
                    16'h265F: data_out = 8'h85;
                    16'h2660: data_out = 8'h86;
                    16'h2661: data_out = 8'h87;
                    16'h2662: data_out = 8'h88;
                    16'h2663: data_out = 8'h89;
                    16'h2664: data_out = 8'h8A;
                    16'h2665: data_out = 8'h8B;
                    16'h2666: data_out = 8'h8C;
                    16'h2667: data_out = 8'h8D;
                    16'h2668: data_out = 8'h8E;
                    16'h2669: data_out = 8'h8F;
                    16'h266A: data_out = 8'h90;
                    16'h266B: data_out = 8'h91;
                    16'h266C: data_out = 8'h92;
                    16'h266D: data_out = 8'h93;
                    16'h266E: data_out = 8'h94;
                    16'h266F: data_out = 8'h95;
                    16'h2670: data_out = 8'h96;
                    16'h2671: data_out = 8'h97;
                    16'h2672: data_out = 8'h98;
                    16'h2673: data_out = 8'h99;
                    16'h2674: data_out = 8'h9A;
                    16'h2675: data_out = 8'h9B;
                    16'h2676: data_out = 8'h9C;
                    16'h2677: data_out = 8'h9D;
                    16'h2678: data_out = 8'h9E;
                    16'h2679: data_out = 8'h9F;
                    16'h267A: data_out = 8'hA0;
                    16'h267B: data_out = 8'hA1;
                    16'h267C: data_out = 8'hA2;
                    16'h267D: data_out = 8'hA3;
                    16'h267E: data_out = 8'hA4;
                    16'h267F: data_out = 8'hA5;
                    16'h2680: data_out = 8'h26;
                    16'h2681: data_out = 8'h25;
                    16'h2682: data_out = 8'h24;
                    16'h2683: data_out = 8'h23;
                    16'h2684: data_out = 8'h22;
                    16'h2685: data_out = 8'h21;
                    16'h2686: data_out = 8'h20;
                    16'h2687: data_out = 8'h1F;
                    16'h2688: data_out = 8'h1E;
                    16'h2689: data_out = 8'h1D;
                    16'h268A: data_out = 8'h1C;
                    16'h268B: data_out = 8'h1B;
                    16'h268C: data_out = 8'h1A;
                    16'h268D: data_out = 8'h19;
                    16'h268E: data_out = 8'h18;
                    16'h268F: data_out = 8'h17;
                    16'h2690: data_out = 8'h16;
                    16'h2691: data_out = 8'h15;
                    16'h2692: data_out = 8'h14;
                    16'h2693: data_out = 8'h13;
                    16'h2694: data_out = 8'h12;
                    16'h2695: data_out = 8'h11;
                    16'h2696: data_out = 8'h10;
                    16'h2697: data_out = 8'hF;
                    16'h2698: data_out = 8'hE;
                    16'h2699: data_out = 8'hD;
                    16'h269A: data_out = 8'hC;
                    16'h269B: data_out = 8'hB;
                    16'h269C: data_out = 8'hA;
                    16'h269D: data_out = 8'h9;
                    16'h269E: data_out = 8'h8;
                    16'h269F: data_out = 8'h7;
                    16'h26A0: data_out = 8'h6;
                    16'h26A1: data_out = 8'h5;
                    16'h26A2: data_out = 8'h4;
                    16'h26A3: data_out = 8'h3;
                    16'h26A4: data_out = 8'h2;
                    16'h26A5: data_out = 8'h1;
                    16'h26A6: data_out = 8'h0;
                    16'h26A7: data_out = 8'h81;
                    16'h26A8: data_out = 8'h82;
                    16'h26A9: data_out = 8'h83;
                    16'h26AA: data_out = 8'h84;
                    16'h26AB: data_out = 8'h85;
                    16'h26AC: data_out = 8'h86;
                    16'h26AD: data_out = 8'h87;
                    16'h26AE: data_out = 8'h88;
                    16'h26AF: data_out = 8'h89;
                    16'h26B0: data_out = 8'h8A;
                    16'h26B1: data_out = 8'h8B;
                    16'h26B2: data_out = 8'h8C;
                    16'h26B3: data_out = 8'h8D;
                    16'h26B4: data_out = 8'h8E;
                    16'h26B5: data_out = 8'h8F;
                    16'h26B6: data_out = 8'h90;
                    16'h26B7: data_out = 8'h91;
                    16'h26B8: data_out = 8'h92;
                    16'h26B9: data_out = 8'h93;
                    16'h26BA: data_out = 8'h94;
                    16'h26BB: data_out = 8'h95;
                    16'h26BC: data_out = 8'h96;
                    16'h26BD: data_out = 8'h97;
                    16'h26BE: data_out = 8'h98;
                    16'h26BF: data_out = 8'h99;
                    16'h26C0: data_out = 8'h9A;
                    16'h26C1: data_out = 8'h9B;
                    16'h26C2: data_out = 8'h9C;
                    16'h26C3: data_out = 8'h9D;
                    16'h26C4: data_out = 8'h9E;
                    16'h26C5: data_out = 8'h9F;
                    16'h26C6: data_out = 8'hA0;
                    16'h26C7: data_out = 8'hA1;
                    16'h26C8: data_out = 8'hA2;
                    16'h26C9: data_out = 8'hA3;
                    16'h26CA: data_out = 8'hA4;
                    16'h26CB: data_out = 8'hA5;
                    16'h26CC: data_out = 8'hA6;
                    16'h26CD: data_out = 8'hA7;
                    16'h26CE: data_out = 8'hA8;
                    16'h26CF: data_out = 8'hA9;
                    16'h26D0: data_out = 8'hAA;
                    16'h26D1: data_out = 8'hAB;
                    16'h26D2: data_out = 8'hAC;
                    16'h26D3: data_out = 8'hAD;
                    16'h26D4: data_out = 8'hAE;
                    16'h26D5: data_out = 8'hAF;
                    16'h26D6: data_out = 8'hB0;
                    16'h26D7: data_out = 8'hB1;
                    16'h26D8: data_out = 8'hB2;
                    16'h26D9: data_out = 8'hB3;
                    16'h26DA: data_out = 8'hB4;
                    16'h26DB: data_out = 8'hB5;
                    16'h26DC: data_out = 8'hB6;
                    16'h26DD: data_out = 8'hB7;
                    16'h26DE: data_out = 8'hB8;
                    16'h26DF: data_out = 8'hB9;
                    16'h26E0: data_out = 8'hBA;
                    16'h26E1: data_out = 8'hBB;
                    16'h26E2: data_out = 8'hBC;
                    16'h26E3: data_out = 8'hBD;
                    16'h26E4: data_out = 8'hBE;
                    16'h26E5: data_out = 8'hBF;
                    16'h26E6: data_out = 8'hC0;
                    16'h26E7: data_out = 8'hC1;
                    16'h26E8: data_out = 8'hC2;
                    16'h26E9: data_out = 8'hC3;
                    16'h26EA: data_out = 8'hC4;
                    16'h26EB: data_out = 8'hC5;
                    16'h26EC: data_out = 8'hC6;
                    16'h26ED: data_out = 8'hC7;
                    16'h26EE: data_out = 8'hC8;
                    16'h26EF: data_out = 8'hC9;
                    16'h26F0: data_out = 8'hCA;
                    16'h26F1: data_out = 8'hCB;
                    16'h26F2: data_out = 8'hCC;
                    16'h26F3: data_out = 8'hCD;
                    16'h26F4: data_out = 8'hCE;
                    16'h26F5: data_out = 8'hCF;
                    16'h26F6: data_out = 8'hD0;
                    16'h26F7: data_out = 8'hD1;
                    16'h26F8: data_out = 8'hD2;
                    16'h26F9: data_out = 8'hD3;
                    16'h26FA: data_out = 8'hD4;
                    16'h26FB: data_out = 8'hD5;
                    16'h26FC: data_out = 8'hD6;
                    16'h26FD: data_out = 8'hD7;
                    16'h26FE: data_out = 8'hD8;
                    16'h26FF: data_out = 8'hD9;
                    16'h2700: data_out = 8'h27;
                    16'h2701: data_out = 8'h28;
                    16'h2702: data_out = 8'h29;
                    16'h2703: data_out = 8'h2A;
                    16'h2704: data_out = 8'h2B;
                    16'h2705: data_out = 8'h2C;
                    16'h2706: data_out = 8'h2D;
                    16'h2707: data_out = 8'h2E;
                    16'h2708: data_out = 8'h2F;
                    16'h2709: data_out = 8'h30;
                    16'h270A: data_out = 8'h31;
                    16'h270B: data_out = 8'h32;
                    16'h270C: data_out = 8'h33;
                    16'h270D: data_out = 8'h34;
                    16'h270E: data_out = 8'h35;
                    16'h270F: data_out = 8'h36;
                    16'h2710: data_out = 8'h37;
                    16'h2711: data_out = 8'h38;
                    16'h2712: data_out = 8'h39;
                    16'h2713: data_out = 8'h3A;
                    16'h2714: data_out = 8'h3B;
                    16'h2715: data_out = 8'h3C;
                    16'h2716: data_out = 8'h3D;
                    16'h2717: data_out = 8'h3E;
                    16'h2718: data_out = 8'h3F;
                    16'h2719: data_out = 8'h40;
                    16'h271A: data_out = 8'h41;
                    16'h271B: data_out = 8'h42;
                    16'h271C: data_out = 8'h43;
                    16'h271D: data_out = 8'h44;
                    16'h271E: data_out = 8'h45;
                    16'h271F: data_out = 8'h46;
                    16'h2720: data_out = 8'h47;
                    16'h2721: data_out = 8'h48;
                    16'h2722: data_out = 8'h49;
                    16'h2723: data_out = 8'h4A;
                    16'h2724: data_out = 8'h4B;
                    16'h2725: data_out = 8'h4C;
                    16'h2726: data_out = 8'h4D;
                    16'h2727: data_out = 8'h4E;
                    16'h2728: data_out = 8'h4F;
                    16'h2729: data_out = 8'h50;
                    16'h272A: data_out = 8'h51;
                    16'h272B: data_out = 8'h52;
                    16'h272C: data_out = 8'h53;
                    16'h272D: data_out = 8'h54;
                    16'h272E: data_out = 8'h55;
                    16'h272F: data_out = 8'h56;
                    16'h2730: data_out = 8'h57;
                    16'h2731: data_out = 8'h58;
                    16'h2732: data_out = 8'h59;
                    16'h2733: data_out = 8'h5A;
                    16'h2734: data_out = 8'h5B;
                    16'h2735: data_out = 8'h5C;
                    16'h2736: data_out = 8'h5D;
                    16'h2737: data_out = 8'h5E;
                    16'h2738: data_out = 8'h5F;
                    16'h2739: data_out = 8'h60;
                    16'h273A: data_out = 8'h61;
                    16'h273B: data_out = 8'h62;
                    16'h273C: data_out = 8'h63;
                    16'h273D: data_out = 8'h64;
                    16'h273E: data_out = 8'h65;
                    16'h273F: data_out = 8'h66;
                    16'h2740: data_out = 8'h67;
                    16'h2741: data_out = 8'h68;
                    16'h2742: data_out = 8'h69;
                    16'h2743: data_out = 8'h6A;
                    16'h2744: data_out = 8'h6B;
                    16'h2745: data_out = 8'h6C;
                    16'h2746: data_out = 8'h6D;
                    16'h2747: data_out = 8'h6E;
                    16'h2748: data_out = 8'h6F;
                    16'h2749: data_out = 8'h70;
                    16'h274A: data_out = 8'h71;
                    16'h274B: data_out = 8'h72;
                    16'h274C: data_out = 8'h73;
                    16'h274D: data_out = 8'h74;
                    16'h274E: data_out = 8'h75;
                    16'h274F: data_out = 8'h76;
                    16'h2750: data_out = 8'h77;
                    16'h2751: data_out = 8'h78;
                    16'h2752: data_out = 8'h79;
                    16'h2753: data_out = 8'h7A;
                    16'h2754: data_out = 8'h7B;
                    16'h2755: data_out = 8'h7C;
                    16'h2756: data_out = 8'h7D;
                    16'h2757: data_out = 8'h7E;
                    16'h2758: data_out = 8'h7F;
                    16'h2759: data_out = 8'h80;
                    16'h275A: data_out = 8'h81;
                    16'h275B: data_out = 8'h82;
                    16'h275C: data_out = 8'h83;
                    16'h275D: data_out = 8'h84;
                    16'h275E: data_out = 8'h85;
                    16'h275F: data_out = 8'h86;
                    16'h2760: data_out = 8'h87;
                    16'h2761: data_out = 8'h88;
                    16'h2762: data_out = 8'h89;
                    16'h2763: data_out = 8'h8A;
                    16'h2764: data_out = 8'h8B;
                    16'h2765: data_out = 8'h8C;
                    16'h2766: data_out = 8'h8D;
                    16'h2767: data_out = 8'h8E;
                    16'h2768: data_out = 8'h8F;
                    16'h2769: data_out = 8'h90;
                    16'h276A: data_out = 8'h91;
                    16'h276B: data_out = 8'h92;
                    16'h276C: data_out = 8'h93;
                    16'h276D: data_out = 8'h94;
                    16'h276E: data_out = 8'h95;
                    16'h276F: data_out = 8'h96;
                    16'h2770: data_out = 8'h97;
                    16'h2771: data_out = 8'h98;
                    16'h2772: data_out = 8'h99;
                    16'h2773: data_out = 8'h9A;
                    16'h2774: data_out = 8'h9B;
                    16'h2775: data_out = 8'h9C;
                    16'h2776: data_out = 8'h9D;
                    16'h2777: data_out = 8'h9E;
                    16'h2778: data_out = 8'h9F;
                    16'h2779: data_out = 8'hA0;
                    16'h277A: data_out = 8'hA1;
                    16'h277B: data_out = 8'hA2;
                    16'h277C: data_out = 8'hA3;
                    16'h277D: data_out = 8'hA4;
                    16'h277E: data_out = 8'hA5;
                    16'h277F: data_out = 8'hA6;
                    16'h2780: data_out = 8'h27;
                    16'h2781: data_out = 8'h26;
                    16'h2782: data_out = 8'h25;
                    16'h2783: data_out = 8'h24;
                    16'h2784: data_out = 8'h23;
                    16'h2785: data_out = 8'h22;
                    16'h2786: data_out = 8'h21;
                    16'h2787: data_out = 8'h20;
                    16'h2788: data_out = 8'h1F;
                    16'h2789: data_out = 8'h1E;
                    16'h278A: data_out = 8'h1D;
                    16'h278B: data_out = 8'h1C;
                    16'h278C: data_out = 8'h1B;
                    16'h278D: data_out = 8'h1A;
                    16'h278E: data_out = 8'h19;
                    16'h278F: data_out = 8'h18;
                    16'h2790: data_out = 8'h17;
                    16'h2791: data_out = 8'h16;
                    16'h2792: data_out = 8'h15;
                    16'h2793: data_out = 8'h14;
                    16'h2794: data_out = 8'h13;
                    16'h2795: data_out = 8'h12;
                    16'h2796: data_out = 8'h11;
                    16'h2797: data_out = 8'h10;
                    16'h2798: data_out = 8'hF;
                    16'h2799: data_out = 8'hE;
                    16'h279A: data_out = 8'hD;
                    16'h279B: data_out = 8'hC;
                    16'h279C: data_out = 8'hB;
                    16'h279D: data_out = 8'hA;
                    16'h279E: data_out = 8'h9;
                    16'h279F: data_out = 8'h8;
                    16'h27A0: data_out = 8'h7;
                    16'h27A1: data_out = 8'h6;
                    16'h27A2: data_out = 8'h5;
                    16'h27A3: data_out = 8'h4;
                    16'h27A4: data_out = 8'h3;
                    16'h27A5: data_out = 8'h2;
                    16'h27A6: data_out = 8'h1;
                    16'h27A7: data_out = 8'h0;
                    16'h27A8: data_out = 8'h81;
                    16'h27A9: data_out = 8'h82;
                    16'h27AA: data_out = 8'h83;
                    16'h27AB: data_out = 8'h84;
                    16'h27AC: data_out = 8'h85;
                    16'h27AD: data_out = 8'h86;
                    16'h27AE: data_out = 8'h87;
                    16'h27AF: data_out = 8'h88;
                    16'h27B0: data_out = 8'h89;
                    16'h27B1: data_out = 8'h8A;
                    16'h27B2: data_out = 8'h8B;
                    16'h27B3: data_out = 8'h8C;
                    16'h27B4: data_out = 8'h8D;
                    16'h27B5: data_out = 8'h8E;
                    16'h27B6: data_out = 8'h8F;
                    16'h27B7: data_out = 8'h90;
                    16'h27B8: data_out = 8'h91;
                    16'h27B9: data_out = 8'h92;
                    16'h27BA: data_out = 8'h93;
                    16'h27BB: data_out = 8'h94;
                    16'h27BC: data_out = 8'h95;
                    16'h27BD: data_out = 8'h96;
                    16'h27BE: data_out = 8'h97;
                    16'h27BF: data_out = 8'h98;
                    16'h27C0: data_out = 8'h99;
                    16'h27C1: data_out = 8'h9A;
                    16'h27C2: data_out = 8'h9B;
                    16'h27C3: data_out = 8'h9C;
                    16'h27C4: data_out = 8'h9D;
                    16'h27C5: data_out = 8'h9E;
                    16'h27C6: data_out = 8'h9F;
                    16'h27C7: data_out = 8'hA0;
                    16'h27C8: data_out = 8'hA1;
                    16'h27C9: data_out = 8'hA2;
                    16'h27CA: data_out = 8'hA3;
                    16'h27CB: data_out = 8'hA4;
                    16'h27CC: data_out = 8'hA5;
                    16'h27CD: data_out = 8'hA6;
                    16'h27CE: data_out = 8'hA7;
                    16'h27CF: data_out = 8'hA8;
                    16'h27D0: data_out = 8'hA9;
                    16'h27D1: data_out = 8'hAA;
                    16'h27D2: data_out = 8'hAB;
                    16'h27D3: data_out = 8'hAC;
                    16'h27D4: data_out = 8'hAD;
                    16'h27D5: data_out = 8'hAE;
                    16'h27D6: data_out = 8'hAF;
                    16'h27D7: data_out = 8'hB0;
                    16'h27D8: data_out = 8'hB1;
                    16'h27D9: data_out = 8'hB2;
                    16'h27DA: data_out = 8'hB3;
                    16'h27DB: data_out = 8'hB4;
                    16'h27DC: data_out = 8'hB5;
                    16'h27DD: data_out = 8'hB6;
                    16'h27DE: data_out = 8'hB7;
                    16'h27DF: data_out = 8'hB8;
                    16'h27E0: data_out = 8'hB9;
                    16'h27E1: data_out = 8'hBA;
                    16'h27E2: data_out = 8'hBB;
                    16'h27E3: data_out = 8'hBC;
                    16'h27E4: data_out = 8'hBD;
                    16'h27E5: data_out = 8'hBE;
                    16'h27E6: data_out = 8'hBF;
                    16'h27E7: data_out = 8'hC0;
                    16'h27E8: data_out = 8'hC1;
                    16'h27E9: data_out = 8'hC2;
                    16'h27EA: data_out = 8'hC3;
                    16'h27EB: data_out = 8'hC4;
                    16'h27EC: data_out = 8'hC5;
                    16'h27ED: data_out = 8'hC6;
                    16'h27EE: data_out = 8'hC7;
                    16'h27EF: data_out = 8'hC8;
                    16'h27F0: data_out = 8'hC9;
                    16'h27F1: data_out = 8'hCA;
                    16'h27F2: data_out = 8'hCB;
                    16'h27F3: data_out = 8'hCC;
                    16'h27F4: data_out = 8'hCD;
                    16'h27F5: data_out = 8'hCE;
                    16'h27F6: data_out = 8'hCF;
                    16'h27F7: data_out = 8'hD0;
                    16'h27F8: data_out = 8'hD1;
                    16'h27F9: data_out = 8'hD2;
                    16'h27FA: data_out = 8'hD3;
                    16'h27FB: data_out = 8'hD4;
                    16'h27FC: data_out = 8'hD5;
                    16'h27FD: data_out = 8'hD6;
                    16'h27FE: data_out = 8'hD7;
                    16'h27FF: data_out = 8'hD8;
                    16'h2800: data_out = 8'h28;
                    16'h2801: data_out = 8'h29;
                    16'h2802: data_out = 8'h2A;
                    16'h2803: data_out = 8'h2B;
                    16'h2804: data_out = 8'h2C;
                    16'h2805: data_out = 8'h2D;
                    16'h2806: data_out = 8'h2E;
                    16'h2807: data_out = 8'h2F;
                    16'h2808: data_out = 8'h30;
                    16'h2809: data_out = 8'h31;
                    16'h280A: data_out = 8'h32;
                    16'h280B: data_out = 8'h33;
                    16'h280C: data_out = 8'h34;
                    16'h280D: data_out = 8'h35;
                    16'h280E: data_out = 8'h36;
                    16'h280F: data_out = 8'h37;
                    16'h2810: data_out = 8'h38;
                    16'h2811: data_out = 8'h39;
                    16'h2812: data_out = 8'h3A;
                    16'h2813: data_out = 8'h3B;
                    16'h2814: data_out = 8'h3C;
                    16'h2815: data_out = 8'h3D;
                    16'h2816: data_out = 8'h3E;
                    16'h2817: data_out = 8'h3F;
                    16'h2818: data_out = 8'h40;
                    16'h2819: data_out = 8'h41;
                    16'h281A: data_out = 8'h42;
                    16'h281B: data_out = 8'h43;
                    16'h281C: data_out = 8'h44;
                    16'h281D: data_out = 8'h45;
                    16'h281E: data_out = 8'h46;
                    16'h281F: data_out = 8'h47;
                    16'h2820: data_out = 8'h48;
                    16'h2821: data_out = 8'h49;
                    16'h2822: data_out = 8'h4A;
                    16'h2823: data_out = 8'h4B;
                    16'h2824: data_out = 8'h4C;
                    16'h2825: data_out = 8'h4D;
                    16'h2826: data_out = 8'h4E;
                    16'h2827: data_out = 8'h4F;
                    16'h2828: data_out = 8'h50;
                    16'h2829: data_out = 8'h51;
                    16'h282A: data_out = 8'h52;
                    16'h282B: data_out = 8'h53;
                    16'h282C: data_out = 8'h54;
                    16'h282D: data_out = 8'h55;
                    16'h282E: data_out = 8'h56;
                    16'h282F: data_out = 8'h57;
                    16'h2830: data_out = 8'h58;
                    16'h2831: data_out = 8'h59;
                    16'h2832: data_out = 8'h5A;
                    16'h2833: data_out = 8'h5B;
                    16'h2834: data_out = 8'h5C;
                    16'h2835: data_out = 8'h5D;
                    16'h2836: data_out = 8'h5E;
                    16'h2837: data_out = 8'h5F;
                    16'h2838: data_out = 8'h60;
                    16'h2839: data_out = 8'h61;
                    16'h283A: data_out = 8'h62;
                    16'h283B: data_out = 8'h63;
                    16'h283C: data_out = 8'h64;
                    16'h283D: data_out = 8'h65;
                    16'h283E: data_out = 8'h66;
                    16'h283F: data_out = 8'h67;
                    16'h2840: data_out = 8'h68;
                    16'h2841: data_out = 8'h69;
                    16'h2842: data_out = 8'h6A;
                    16'h2843: data_out = 8'h6B;
                    16'h2844: data_out = 8'h6C;
                    16'h2845: data_out = 8'h6D;
                    16'h2846: data_out = 8'h6E;
                    16'h2847: data_out = 8'h6F;
                    16'h2848: data_out = 8'h70;
                    16'h2849: data_out = 8'h71;
                    16'h284A: data_out = 8'h72;
                    16'h284B: data_out = 8'h73;
                    16'h284C: data_out = 8'h74;
                    16'h284D: data_out = 8'h75;
                    16'h284E: data_out = 8'h76;
                    16'h284F: data_out = 8'h77;
                    16'h2850: data_out = 8'h78;
                    16'h2851: data_out = 8'h79;
                    16'h2852: data_out = 8'h7A;
                    16'h2853: data_out = 8'h7B;
                    16'h2854: data_out = 8'h7C;
                    16'h2855: data_out = 8'h7D;
                    16'h2856: data_out = 8'h7E;
                    16'h2857: data_out = 8'h7F;
                    16'h2858: data_out = 8'h80;
                    16'h2859: data_out = 8'h81;
                    16'h285A: data_out = 8'h82;
                    16'h285B: data_out = 8'h83;
                    16'h285C: data_out = 8'h84;
                    16'h285D: data_out = 8'h85;
                    16'h285E: data_out = 8'h86;
                    16'h285F: data_out = 8'h87;
                    16'h2860: data_out = 8'h88;
                    16'h2861: data_out = 8'h89;
                    16'h2862: data_out = 8'h8A;
                    16'h2863: data_out = 8'h8B;
                    16'h2864: data_out = 8'h8C;
                    16'h2865: data_out = 8'h8D;
                    16'h2866: data_out = 8'h8E;
                    16'h2867: data_out = 8'h8F;
                    16'h2868: data_out = 8'h90;
                    16'h2869: data_out = 8'h91;
                    16'h286A: data_out = 8'h92;
                    16'h286B: data_out = 8'h93;
                    16'h286C: data_out = 8'h94;
                    16'h286D: data_out = 8'h95;
                    16'h286E: data_out = 8'h96;
                    16'h286F: data_out = 8'h97;
                    16'h2870: data_out = 8'h98;
                    16'h2871: data_out = 8'h99;
                    16'h2872: data_out = 8'h9A;
                    16'h2873: data_out = 8'h9B;
                    16'h2874: data_out = 8'h9C;
                    16'h2875: data_out = 8'h9D;
                    16'h2876: data_out = 8'h9E;
                    16'h2877: data_out = 8'h9F;
                    16'h2878: data_out = 8'hA0;
                    16'h2879: data_out = 8'hA1;
                    16'h287A: data_out = 8'hA2;
                    16'h287B: data_out = 8'hA3;
                    16'h287C: data_out = 8'hA4;
                    16'h287D: data_out = 8'hA5;
                    16'h287E: data_out = 8'hA6;
                    16'h287F: data_out = 8'hA7;
                    16'h2880: data_out = 8'h28;
                    16'h2881: data_out = 8'h27;
                    16'h2882: data_out = 8'h26;
                    16'h2883: data_out = 8'h25;
                    16'h2884: data_out = 8'h24;
                    16'h2885: data_out = 8'h23;
                    16'h2886: data_out = 8'h22;
                    16'h2887: data_out = 8'h21;
                    16'h2888: data_out = 8'h20;
                    16'h2889: data_out = 8'h1F;
                    16'h288A: data_out = 8'h1E;
                    16'h288B: data_out = 8'h1D;
                    16'h288C: data_out = 8'h1C;
                    16'h288D: data_out = 8'h1B;
                    16'h288E: data_out = 8'h1A;
                    16'h288F: data_out = 8'h19;
                    16'h2890: data_out = 8'h18;
                    16'h2891: data_out = 8'h17;
                    16'h2892: data_out = 8'h16;
                    16'h2893: data_out = 8'h15;
                    16'h2894: data_out = 8'h14;
                    16'h2895: data_out = 8'h13;
                    16'h2896: data_out = 8'h12;
                    16'h2897: data_out = 8'h11;
                    16'h2898: data_out = 8'h10;
                    16'h2899: data_out = 8'hF;
                    16'h289A: data_out = 8'hE;
                    16'h289B: data_out = 8'hD;
                    16'h289C: data_out = 8'hC;
                    16'h289D: data_out = 8'hB;
                    16'h289E: data_out = 8'hA;
                    16'h289F: data_out = 8'h9;
                    16'h28A0: data_out = 8'h8;
                    16'h28A1: data_out = 8'h7;
                    16'h28A2: data_out = 8'h6;
                    16'h28A3: data_out = 8'h5;
                    16'h28A4: data_out = 8'h4;
                    16'h28A5: data_out = 8'h3;
                    16'h28A6: data_out = 8'h2;
                    16'h28A7: data_out = 8'h1;
                    16'h28A8: data_out = 8'h0;
                    16'h28A9: data_out = 8'h81;
                    16'h28AA: data_out = 8'h82;
                    16'h28AB: data_out = 8'h83;
                    16'h28AC: data_out = 8'h84;
                    16'h28AD: data_out = 8'h85;
                    16'h28AE: data_out = 8'h86;
                    16'h28AF: data_out = 8'h87;
                    16'h28B0: data_out = 8'h88;
                    16'h28B1: data_out = 8'h89;
                    16'h28B2: data_out = 8'h8A;
                    16'h28B3: data_out = 8'h8B;
                    16'h28B4: data_out = 8'h8C;
                    16'h28B5: data_out = 8'h8D;
                    16'h28B6: data_out = 8'h8E;
                    16'h28B7: data_out = 8'h8F;
                    16'h28B8: data_out = 8'h90;
                    16'h28B9: data_out = 8'h91;
                    16'h28BA: data_out = 8'h92;
                    16'h28BB: data_out = 8'h93;
                    16'h28BC: data_out = 8'h94;
                    16'h28BD: data_out = 8'h95;
                    16'h28BE: data_out = 8'h96;
                    16'h28BF: data_out = 8'h97;
                    16'h28C0: data_out = 8'h98;
                    16'h28C1: data_out = 8'h99;
                    16'h28C2: data_out = 8'h9A;
                    16'h28C3: data_out = 8'h9B;
                    16'h28C4: data_out = 8'h9C;
                    16'h28C5: data_out = 8'h9D;
                    16'h28C6: data_out = 8'h9E;
                    16'h28C7: data_out = 8'h9F;
                    16'h28C8: data_out = 8'hA0;
                    16'h28C9: data_out = 8'hA1;
                    16'h28CA: data_out = 8'hA2;
                    16'h28CB: data_out = 8'hA3;
                    16'h28CC: data_out = 8'hA4;
                    16'h28CD: data_out = 8'hA5;
                    16'h28CE: data_out = 8'hA6;
                    16'h28CF: data_out = 8'hA7;
                    16'h28D0: data_out = 8'hA8;
                    16'h28D1: data_out = 8'hA9;
                    16'h28D2: data_out = 8'hAA;
                    16'h28D3: data_out = 8'hAB;
                    16'h28D4: data_out = 8'hAC;
                    16'h28D5: data_out = 8'hAD;
                    16'h28D6: data_out = 8'hAE;
                    16'h28D7: data_out = 8'hAF;
                    16'h28D8: data_out = 8'hB0;
                    16'h28D9: data_out = 8'hB1;
                    16'h28DA: data_out = 8'hB2;
                    16'h28DB: data_out = 8'hB3;
                    16'h28DC: data_out = 8'hB4;
                    16'h28DD: data_out = 8'hB5;
                    16'h28DE: data_out = 8'hB6;
                    16'h28DF: data_out = 8'hB7;
                    16'h28E0: data_out = 8'hB8;
                    16'h28E1: data_out = 8'hB9;
                    16'h28E2: data_out = 8'hBA;
                    16'h28E3: data_out = 8'hBB;
                    16'h28E4: data_out = 8'hBC;
                    16'h28E5: data_out = 8'hBD;
                    16'h28E6: data_out = 8'hBE;
                    16'h28E7: data_out = 8'hBF;
                    16'h28E8: data_out = 8'hC0;
                    16'h28E9: data_out = 8'hC1;
                    16'h28EA: data_out = 8'hC2;
                    16'h28EB: data_out = 8'hC3;
                    16'h28EC: data_out = 8'hC4;
                    16'h28ED: data_out = 8'hC5;
                    16'h28EE: data_out = 8'hC6;
                    16'h28EF: data_out = 8'hC7;
                    16'h28F0: data_out = 8'hC8;
                    16'h28F1: data_out = 8'hC9;
                    16'h28F2: data_out = 8'hCA;
                    16'h28F3: data_out = 8'hCB;
                    16'h28F4: data_out = 8'hCC;
                    16'h28F5: data_out = 8'hCD;
                    16'h28F6: data_out = 8'hCE;
                    16'h28F7: data_out = 8'hCF;
                    16'h28F8: data_out = 8'hD0;
                    16'h28F9: data_out = 8'hD1;
                    16'h28FA: data_out = 8'hD2;
                    16'h28FB: data_out = 8'hD3;
                    16'h28FC: data_out = 8'hD4;
                    16'h28FD: data_out = 8'hD5;
                    16'h28FE: data_out = 8'hD6;
                    16'h28FF: data_out = 8'hD7;
                    16'h2900: data_out = 8'h29;
                    16'h2901: data_out = 8'h2A;
                    16'h2902: data_out = 8'h2B;
                    16'h2903: data_out = 8'h2C;
                    16'h2904: data_out = 8'h2D;
                    16'h2905: data_out = 8'h2E;
                    16'h2906: data_out = 8'h2F;
                    16'h2907: data_out = 8'h30;
                    16'h2908: data_out = 8'h31;
                    16'h2909: data_out = 8'h32;
                    16'h290A: data_out = 8'h33;
                    16'h290B: data_out = 8'h34;
                    16'h290C: data_out = 8'h35;
                    16'h290D: data_out = 8'h36;
                    16'h290E: data_out = 8'h37;
                    16'h290F: data_out = 8'h38;
                    16'h2910: data_out = 8'h39;
                    16'h2911: data_out = 8'h3A;
                    16'h2912: data_out = 8'h3B;
                    16'h2913: data_out = 8'h3C;
                    16'h2914: data_out = 8'h3D;
                    16'h2915: data_out = 8'h3E;
                    16'h2916: data_out = 8'h3F;
                    16'h2917: data_out = 8'h40;
                    16'h2918: data_out = 8'h41;
                    16'h2919: data_out = 8'h42;
                    16'h291A: data_out = 8'h43;
                    16'h291B: data_out = 8'h44;
                    16'h291C: data_out = 8'h45;
                    16'h291D: data_out = 8'h46;
                    16'h291E: data_out = 8'h47;
                    16'h291F: data_out = 8'h48;
                    16'h2920: data_out = 8'h49;
                    16'h2921: data_out = 8'h4A;
                    16'h2922: data_out = 8'h4B;
                    16'h2923: data_out = 8'h4C;
                    16'h2924: data_out = 8'h4D;
                    16'h2925: data_out = 8'h4E;
                    16'h2926: data_out = 8'h4F;
                    16'h2927: data_out = 8'h50;
                    16'h2928: data_out = 8'h51;
                    16'h2929: data_out = 8'h52;
                    16'h292A: data_out = 8'h53;
                    16'h292B: data_out = 8'h54;
                    16'h292C: data_out = 8'h55;
                    16'h292D: data_out = 8'h56;
                    16'h292E: data_out = 8'h57;
                    16'h292F: data_out = 8'h58;
                    16'h2930: data_out = 8'h59;
                    16'h2931: data_out = 8'h5A;
                    16'h2932: data_out = 8'h5B;
                    16'h2933: data_out = 8'h5C;
                    16'h2934: data_out = 8'h5D;
                    16'h2935: data_out = 8'h5E;
                    16'h2936: data_out = 8'h5F;
                    16'h2937: data_out = 8'h60;
                    16'h2938: data_out = 8'h61;
                    16'h2939: data_out = 8'h62;
                    16'h293A: data_out = 8'h63;
                    16'h293B: data_out = 8'h64;
                    16'h293C: data_out = 8'h65;
                    16'h293D: data_out = 8'h66;
                    16'h293E: data_out = 8'h67;
                    16'h293F: data_out = 8'h68;
                    16'h2940: data_out = 8'h69;
                    16'h2941: data_out = 8'h6A;
                    16'h2942: data_out = 8'h6B;
                    16'h2943: data_out = 8'h6C;
                    16'h2944: data_out = 8'h6D;
                    16'h2945: data_out = 8'h6E;
                    16'h2946: data_out = 8'h6F;
                    16'h2947: data_out = 8'h70;
                    16'h2948: data_out = 8'h71;
                    16'h2949: data_out = 8'h72;
                    16'h294A: data_out = 8'h73;
                    16'h294B: data_out = 8'h74;
                    16'h294C: data_out = 8'h75;
                    16'h294D: data_out = 8'h76;
                    16'h294E: data_out = 8'h77;
                    16'h294F: data_out = 8'h78;
                    16'h2950: data_out = 8'h79;
                    16'h2951: data_out = 8'h7A;
                    16'h2952: data_out = 8'h7B;
                    16'h2953: data_out = 8'h7C;
                    16'h2954: data_out = 8'h7D;
                    16'h2955: data_out = 8'h7E;
                    16'h2956: data_out = 8'h7F;
                    16'h2957: data_out = 8'h80;
                    16'h2958: data_out = 8'h81;
                    16'h2959: data_out = 8'h82;
                    16'h295A: data_out = 8'h83;
                    16'h295B: data_out = 8'h84;
                    16'h295C: data_out = 8'h85;
                    16'h295D: data_out = 8'h86;
                    16'h295E: data_out = 8'h87;
                    16'h295F: data_out = 8'h88;
                    16'h2960: data_out = 8'h89;
                    16'h2961: data_out = 8'h8A;
                    16'h2962: data_out = 8'h8B;
                    16'h2963: data_out = 8'h8C;
                    16'h2964: data_out = 8'h8D;
                    16'h2965: data_out = 8'h8E;
                    16'h2966: data_out = 8'h8F;
                    16'h2967: data_out = 8'h90;
                    16'h2968: data_out = 8'h91;
                    16'h2969: data_out = 8'h92;
                    16'h296A: data_out = 8'h93;
                    16'h296B: data_out = 8'h94;
                    16'h296C: data_out = 8'h95;
                    16'h296D: data_out = 8'h96;
                    16'h296E: data_out = 8'h97;
                    16'h296F: data_out = 8'h98;
                    16'h2970: data_out = 8'h99;
                    16'h2971: data_out = 8'h9A;
                    16'h2972: data_out = 8'h9B;
                    16'h2973: data_out = 8'h9C;
                    16'h2974: data_out = 8'h9D;
                    16'h2975: data_out = 8'h9E;
                    16'h2976: data_out = 8'h9F;
                    16'h2977: data_out = 8'hA0;
                    16'h2978: data_out = 8'hA1;
                    16'h2979: data_out = 8'hA2;
                    16'h297A: data_out = 8'hA3;
                    16'h297B: data_out = 8'hA4;
                    16'h297C: data_out = 8'hA5;
                    16'h297D: data_out = 8'hA6;
                    16'h297E: data_out = 8'hA7;
                    16'h297F: data_out = 8'hA8;
                    16'h2980: data_out = 8'h29;
                    16'h2981: data_out = 8'h28;
                    16'h2982: data_out = 8'h27;
                    16'h2983: data_out = 8'h26;
                    16'h2984: data_out = 8'h25;
                    16'h2985: data_out = 8'h24;
                    16'h2986: data_out = 8'h23;
                    16'h2987: data_out = 8'h22;
                    16'h2988: data_out = 8'h21;
                    16'h2989: data_out = 8'h20;
                    16'h298A: data_out = 8'h1F;
                    16'h298B: data_out = 8'h1E;
                    16'h298C: data_out = 8'h1D;
                    16'h298D: data_out = 8'h1C;
                    16'h298E: data_out = 8'h1B;
                    16'h298F: data_out = 8'h1A;
                    16'h2990: data_out = 8'h19;
                    16'h2991: data_out = 8'h18;
                    16'h2992: data_out = 8'h17;
                    16'h2993: data_out = 8'h16;
                    16'h2994: data_out = 8'h15;
                    16'h2995: data_out = 8'h14;
                    16'h2996: data_out = 8'h13;
                    16'h2997: data_out = 8'h12;
                    16'h2998: data_out = 8'h11;
                    16'h2999: data_out = 8'h10;
                    16'h299A: data_out = 8'hF;
                    16'h299B: data_out = 8'hE;
                    16'h299C: data_out = 8'hD;
                    16'h299D: data_out = 8'hC;
                    16'h299E: data_out = 8'hB;
                    16'h299F: data_out = 8'hA;
                    16'h29A0: data_out = 8'h9;
                    16'h29A1: data_out = 8'h8;
                    16'h29A2: data_out = 8'h7;
                    16'h29A3: data_out = 8'h6;
                    16'h29A4: data_out = 8'h5;
                    16'h29A5: data_out = 8'h4;
                    16'h29A6: data_out = 8'h3;
                    16'h29A7: data_out = 8'h2;
                    16'h29A8: data_out = 8'h1;
                    16'h29A9: data_out = 8'h0;
                    16'h29AA: data_out = 8'h81;
                    16'h29AB: data_out = 8'h82;
                    16'h29AC: data_out = 8'h83;
                    16'h29AD: data_out = 8'h84;
                    16'h29AE: data_out = 8'h85;
                    16'h29AF: data_out = 8'h86;
                    16'h29B0: data_out = 8'h87;
                    16'h29B1: data_out = 8'h88;
                    16'h29B2: data_out = 8'h89;
                    16'h29B3: data_out = 8'h8A;
                    16'h29B4: data_out = 8'h8B;
                    16'h29B5: data_out = 8'h8C;
                    16'h29B6: data_out = 8'h8D;
                    16'h29B7: data_out = 8'h8E;
                    16'h29B8: data_out = 8'h8F;
                    16'h29B9: data_out = 8'h90;
                    16'h29BA: data_out = 8'h91;
                    16'h29BB: data_out = 8'h92;
                    16'h29BC: data_out = 8'h93;
                    16'h29BD: data_out = 8'h94;
                    16'h29BE: data_out = 8'h95;
                    16'h29BF: data_out = 8'h96;
                    16'h29C0: data_out = 8'h97;
                    16'h29C1: data_out = 8'h98;
                    16'h29C2: data_out = 8'h99;
                    16'h29C3: data_out = 8'h9A;
                    16'h29C4: data_out = 8'h9B;
                    16'h29C5: data_out = 8'h9C;
                    16'h29C6: data_out = 8'h9D;
                    16'h29C7: data_out = 8'h9E;
                    16'h29C8: data_out = 8'h9F;
                    16'h29C9: data_out = 8'hA0;
                    16'h29CA: data_out = 8'hA1;
                    16'h29CB: data_out = 8'hA2;
                    16'h29CC: data_out = 8'hA3;
                    16'h29CD: data_out = 8'hA4;
                    16'h29CE: data_out = 8'hA5;
                    16'h29CF: data_out = 8'hA6;
                    16'h29D0: data_out = 8'hA7;
                    16'h29D1: data_out = 8'hA8;
                    16'h29D2: data_out = 8'hA9;
                    16'h29D3: data_out = 8'hAA;
                    16'h29D4: data_out = 8'hAB;
                    16'h29D5: data_out = 8'hAC;
                    16'h29D6: data_out = 8'hAD;
                    16'h29D7: data_out = 8'hAE;
                    16'h29D8: data_out = 8'hAF;
                    16'h29D9: data_out = 8'hB0;
                    16'h29DA: data_out = 8'hB1;
                    16'h29DB: data_out = 8'hB2;
                    16'h29DC: data_out = 8'hB3;
                    16'h29DD: data_out = 8'hB4;
                    16'h29DE: data_out = 8'hB5;
                    16'h29DF: data_out = 8'hB6;
                    16'h29E0: data_out = 8'hB7;
                    16'h29E1: data_out = 8'hB8;
                    16'h29E2: data_out = 8'hB9;
                    16'h29E3: data_out = 8'hBA;
                    16'h29E4: data_out = 8'hBB;
                    16'h29E5: data_out = 8'hBC;
                    16'h29E6: data_out = 8'hBD;
                    16'h29E7: data_out = 8'hBE;
                    16'h29E8: data_out = 8'hBF;
                    16'h29E9: data_out = 8'hC0;
                    16'h29EA: data_out = 8'hC1;
                    16'h29EB: data_out = 8'hC2;
                    16'h29EC: data_out = 8'hC3;
                    16'h29ED: data_out = 8'hC4;
                    16'h29EE: data_out = 8'hC5;
                    16'h29EF: data_out = 8'hC6;
                    16'h29F0: data_out = 8'hC7;
                    16'h29F1: data_out = 8'hC8;
                    16'h29F2: data_out = 8'hC9;
                    16'h29F3: data_out = 8'hCA;
                    16'h29F4: data_out = 8'hCB;
                    16'h29F5: data_out = 8'hCC;
                    16'h29F6: data_out = 8'hCD;
                    16'h29F7: data_out = 8'hCE;
                    16'h29F8: data_out = 8'hCF;
                    16'h29F9: data_out = 8'hD0;
                    16'h29FA: data_out = 8'hD1;
                    16'h29FB: data_out = 8'hD2;
                    16'h29FC: data_out = 8'hD3;
                    16'h29FD: data_out = 8'hD4;
                    16'h29FE: data_out = 8'hD5;
                    16'h29FF: data_out = 8'hD6;
                    16'h2A00: data_out = 8'h2A;
                    16'h2A01: data_out = 8'h2B;
                    16'h2A02: data_out = 8'h2C;
                    16'h2A03: data_out = 8'h2D;
                    16'h2A04: data_out = 8'h2E;
                    16'h2A05: data_out = 8'h2F;
                    16'h2A06: data_out = 8'h30;
                    16'h2A07: data_out = 8'h31;
                    16'h2A08: data_out = 8'h32;
                    16'h2A09: data_out = 8'h33;
                    16'h2A0A: data_out = 8'h34;
                    16'h2A0B: data_out = 8'h35;
                    16'h2A0C: data_out = 8'h36;
                    16'h2A0D: data_out = 8'h37;
                    16'h2A0E: data_out = 8'h38;
                    16'h2A0F: data_out = 8'h39;
                    16'h2A10: data_out = 8'h3A;
                    16'h2A11: data_out = 8'h3B;
                    16'h2A12: data_out = 8'h3C;
                    16'h2A13: data_out = 8'h3D;
                    16'h2A14: data_out = 8'h3E;
                    16'h2A15: data_out = 8'h3F;
                    16'h2A16: data_out = 8'h40;
                    16'h2A17: data_out = 8'h41;
                    16'h2A18: data_out = 8'h42;
                    16'h2A19: data_out = 8'h43;
                    16'h2A1A: data_out = 8'h44;
                    16'h2A1B: data_out = 8'h45;
                    16'h2A1C: data_out = 8'h46;
                    16'h2A1D: data_out = 8'h47;
                    16'h2A1E: data_out = 8'h48;
                    16'h2A1F: data_out = 8'h49;
                    16'h2A20: data_out = 8'h4A;
                    16'h2A21: data_out = 8'h4B;
                    16'h2A22: data_out = 8'h4C;
                    16'h2A23: data_out = 8'h4D;
                    16'h2A24: data_out = 8'h4E;
                    16'h2A25: data_out = 8'h4F;
                    16'h2A26: data_out = 8'h50;
                    16'h2A27: data_out = 8'h51;
                    16'h2A28: data_out = 8'h52;
                    16'h2A29: data_out = 8'h53;
                    16'h2A2A: data_out = 8'h54;
                    16'h2A2B: data_out = 8'h55;
                    16'h2A2C: data_out = 8'h56;
                    16'h2A2D: data_out = 8'h57;
                    16'h2A2E: data_out = 8'h58;
                    16'h2A2F: data_out = 8'h59;
                    16'h2A30: data_out = 8'h5A;
                    16'h2A31: data_out = 8'h5B;
                    16'h2A32: data_out = 8'h5C;
                    16'h2A33: data_out = 8'h5D;
                    16'h2A34: data_out = 8'h5E;
                    16'h2A35: data_out = 8'h5F;
                    16'h2A36: data_out = 8'h60;
                    16'h2A37: data_out = 8'h61;
                    16'h2A38: data_out = 8'h62;
                    16'h2A39: data_out = 8'h63;
                    16'h2A3A: data_out = 8'h64;
                    16'h2A3B: data_out = 8'h65;
                    16'h2A3C: data_out = 8'h66;
                    16'h2A3D: data_out = 8'h67;
                    16'h2A3E: data_out = 8'h68;
                    16'h2A3F: data_out = 8'h69;
                    16'h2A40: data_out = 8'h6A;
                    16'h2A41: data_out = 8'h6B;
                    16'h2A42: data_out = 8'h6C;
                    16'h2A43: data_out = 8'h6D;
                    16'h2A44: data_out = 8'h6E;
                    16'h2A45: data_out = 8'h6F;
                    16'h2A46: data_out = 8'h70;
                    16'h2A47: data_out = 8'h71;
                    16'h2A48: data_out = 8'h72;
                    16'h2A49: data_out = 8'h73;
                    16'h2A4A: data_out = 8'h74;
                    16'h2A4B: data_out = 8'h75;
                    16'h2A4C: data_out = 8'h76;
                    16'h2A4D: data_out = 8'h77;
                    16'h2A4E: data_out = 8'h78;
                    16'h2A4F: data_out = 8'h79;
                    16'h2A50: data_out = 8'h7A;
                    16'h2A51: data_out = 8'h7B;
                    16'h2A52: data_out = 8'h7C;
                    16'h2A53: data_out = 8'h7D;
                    16'h2A54: data_out = 8'h7E;
                    16'h2A55: data_out = 8'h7F;
                    16'h2A56: data_out = 8'h80;
                    16'h2A57: data_out = 8'h81;
                    16'h2A58: data_out = 8'h82;
                    16'h2A59: data_out = 8'h83;
                    16'h2A5A: data_out = 8'h84;
                    16'h2A5B: data_out = 8'h85;
                    16'h2A5C: data_out = 8'h86;
                    16'h2A5D: data_out = 8'h87;
                    16'h2A5E: data_out = 8'h88;
                    16'h2A5F: data_out = 8'h89;
                    16'h2A60: data_out = 8'h8A;
                    16'h2A61: data_out = 8'h8B;
                    16'h2A62: data_out = 8'h8C;
                    16'h2A63: data_out = 8'h8D;
                    16'h2A64: data_out = 8'h8E;
                    16'h2A65: data_out = 8'h8F;
                    16'h2A66: data_out = 8'h90;
                    16'h2A67: data_out = 8'h91;
                    16'h2A68: data_out = 8'h92;
                    16'h2A69: data_out = 8'h93;
                    16'h2A6A: data_out = 8'h94;
                    16'h2A6B: data_out = 8'h95;
                    16'h2A6C: data_out = 8'h96;
                    16'h2A6D: data_out = 8'h97;
                    16'h2A6E: data_out = 8'h98;
                    16'h2A6F: data_out = 8'h99;
                    16'h2A70: data_out = 8'h9A;
                    16'h2A71: data_out = 8'h9B;
                    16'h2A72: data_out = 8'h9C;
                    16'h2A73: data_out = 8'h9D;
                    16'h2A74: data_out = 8'h9E;
                    16'h2A75: data_out = 8'h9F;
                    16'h2A76: data_out = 8'hA0;
                    16'h2A77: data_out = 8'hA1;
                    16'h2A78: data_out = 8'hA2;
                    16'h2A79: data_out = 8'hA3;
                    16'h2A7A: data_out = 8'hA4;
                    16'h2A7B: data_out = 8'hA5;
                    16'h2A7C: data_out = 8'hA6;
                    16'h2A7D: data_out = 8'hA7;
                    16'h2A7E: data_out = 8'hA8;
                    16'h2A7F: data_out = 8'hA9;
                    16'h2A80: data_out = 8'h2A;
                    16'h2A81: data_out = 8'h29;
                    16'h2A82: data_out = 8'h28;
                    16'h2A83: data_out = 8'h27;
                    16'h2A84: data_out = 8'h26;
                    16'h2A85: data_out = 8'h25;
                    16'h2A86: data_out = 8'h24;
                    16'h2A87: data_out = 8'h23;
                    16'h2A88: data_out = 8'h22;
                    16'h2A89: data_out = 8'h21;
                    16'h2A8A: data_out = 8'h20;
                    16'h2A8B: data_out = 8'h1F;
                    16'h2A8C: data_out = 8'h1E;
                    16'h2A8D: data_out = 8'h1D;
                    16'h2A8E: data_out = 8'h1C;
                    16'h2A8F: data_out = 8'h1B;
                    16'h2A90: data_out = 8'h1A;
                    16'h2A91: data_out = 8'h19;
                    16'h2A92: data_out = 8'h18;
                    16'h2A93: data_out = 8'h17;
                    16'h2A94: data_out = 8'h16;
                    16'h2A95: data_out = 8'h15;
                    16'h2A96: data_out = 8'h14;
                    16'h2A97: data_out = 8'h13;
                    16'h2A98: data_out = 8'h12;
                    16'h2A99: data_out = 8'h11;
                    16'h2A9A: data_out = 8'h10;
                    16'h2A9B: data_out = 8'hF;
                    16'h2A9C: data_out = 8'hE;
                    16'h2A9D: data_out = 8'hD;
                    16'h2A9E: data_out = 8'hC;
                    16'h2A9F: data_out = 8'hB;
                    16'h2AA0: data_out = 8'hA;
                    16'h2AA1: data_out = 8'h9;
                    16'h2AA2: data_out = 8'h8;
                    16'h2AA3: data_out = 8'h7;
                    16'h2AA4: data_out = 8'h6;
                    16'h2AA5: data_out = 8'h5;
                    16'h2AA6: data_out = 8'h4;
                    16'h2AA7: data_out = 8'h3;
                    16'h2AA8: data_out = 8'h2;
                    16'h2AA9: data_out = 8'h1;
                    16'h2AAA: data_out = 8'h0;
                    16'h2AAB: data_out = 8'h81;
                    16'h2AAC: data_out = 8'h82;
                    16'h2AAD: data_out = 8'h83;
                    16'h2AAE: data_out = 8'h84;
                    16'h2AAF: data_out = 8'h85;
                    16'h2AB0: data_out = 8'h86;
                    16'h2AB1: data_out = 8'h87;
                    16'h2AB2: data_out = 8'h88;
                    16'h2AB3: data_out = 8'h89;
                    16'h2AB4: data_out = 8'h8A;
                    16'h2AB5: data_out = 8'h8B;
                    16'h2AB6: data_out = 8'h8C;
                    16'h2AB7: data_out = 8'h8D;
                    16'h2AB8: data_out = 8'h8E;
                    16'h2AB9: data_out = 8'h8F;
                    16'h2ABA: data_out = 8'h90;
                    16'h2ABB: data_out = 8'h91;
                    16'h2ABC: data_out = 8'h92;
                    16'h2ABD: data_out = 8'h93;
                    16'h2ABE: data_out = 8'h94;
                    16'h2ABF: data_out = 8'h95;
                    16'h2AC0: data_out = 8'h96;
                    16'h2AC1: data_out = 8'h97;
                    16'h2AC2: data_out = 8'h98;
                    16'h2AC3: data_out = 8'h99;
                    16'h2AC4: data_out = 8'h9A;
                    16'h2AC5: data_out = 8'h9B;
                    16'h2AC6: data_out = 8'h9C;
                    16'h2AC7: data_out = 8'h9D;
                    16'h2AC8: data_out = 8'h9E;
                    16'h2AC9: data_out = 8'h9F;
                    16'h2ACA: data_out = 8'hA0;
                    16'h2ACB: data_out = 8'hA1;
                    16'h2ACC: data_out = 8'hA2;
                    16'h2ACD: data_out = 8'hA3;
                    16'h2ACE: data_out = 8'hA4;
                    16'h2ACF: data_out = 8'hA5;
                    16'h2AD0: data_out = 8'hA6;
                    16'h2AD1: data_out = 8'hA7;
                    16'h2AD2: data_out = 8'hA8;
                    16'h2AD3: data_out = 8'hA9;
                    16'h2AD4: data_out = 8'hAA;
                    16'h2AD5: data_out = 8'hAB;
                    16'h2AD6: data_out = 8'hAC;
                    16'h2AD7: data_out = 8'hAD;
                    16'h2AD8: data_out = 8'hAE;
                    16'h2AD9: data_out = 8'hAF;
                    16'h2ADA: data_out = 8'hB0;
                    16'h2ADB: data_out = 8'hB1;
                    16'h2ADC: data_out = 8'hB2;
                    16'h2ADD: data_out = 8'hB3;
                    16'h2ADE: data_out = 8'hB4;
                    16'h2ADF: data_out = 8'hB5;
                    16'h2AE0: data_out = 8'hB6;
                    16'h2AE1: data_out = 8'hB7;
                    16'h2AE2: data_out = 8'hB8;
                    16'h2AE3: data_out = 8'hB9;
                    16'h2AE4: data_out = 8'hBA;
                    16'h2AE5: data_out = 8'hBB;
                    16'h2AE6: data_out = 8'hBC;
                    16'h2AE7: data_out = 8'hBD;
                    16'h2AE8: data_out = 8'hBE;
                    16'h2AE9: data_out = 8'hBF;
                    16'h2AEA: data_out = 8'hC0;
                    16'h2AEB: data_out = 8'hC1;
                    16'h2AEC: data_out = 8'hC2;
                    16'h2AED: data_out = 8'hC3;
                    16'h2AEE: data_out = 8'hC4;
                    16'h2AEF: data_out = 8'hC5;
                    16'h2AF0: data_out = 8'hC6;
                    16'h2AF1: data_out = 8'hC7;
                    16'h2AF2: data_out = 8'hC8;
                    16'h2AF3: data_out = 8'hC9;
                    16'h2AF4: data_out = 8'hCA;
                    16'h2AF5: data_out = 8'hCB;
                    16'h2AF6: data_out = 8'hCC;
                    16'h2AF7: data_out = 8'hCD;
                    16'h2AF8: data_out = 8'hCE;
                    16'h2AF9: data_out = 8'hCF;
                    16'h2AFA: data_out = 8'hD0;
                    16'h2AFB: data_out = 8'hD1;
                    16'h2AFC: data_out = 8'hD2;
                    16'h2AFD: data_out = 8'hD3;
                    16'h2AFE: data_out = 8'hD4;
                    16'h2AFF: data_out = 8'hD5;
                    16'h2B00: data_out = 8'h2B;
                    16'h2B01: data_out = 8'h2C;
                    16'h2B02: data_out = 8'h2D;
                    16'h2B03: data_out = 8'h2E;
                    16'h2B04: data_out = 8'h2F;
                    16'h2B05: data_out = 8'h30;
                    16'h2B06: data_out = 8'h31;
                    16'h2B07: data_out = 8'h32;
                    16'h2B08: data_out = 8'h33;
                    16'h2B09: data_out = 8'h34;
                    16'h2B0A: data_out = 8'h35;
                    16'h2B0B: data_out = 8'h36;
                    16'h2B0C: data_out = 8'h37;
                    16'h2B0D: data_out = 8'h38;
                    16'h2B0E: data_out = 8'h39;
                    16'h2B0F: data_out = 8'h3A;
                    16'h2B10: data_out = 8'h3B;
                    16'h2B11: data_out = 8'h3C;
                    16'h2B12: data_out = 8'h3D;
                    16'h2B13: data_out = 8'h3E;
                    16'h2B14: data_out = 8'h3F;
                    16'h2B15: data_out = 8'h40;
                    16'h2B16: data_out = 8'h41;
                    16'h2B17: data_out = 8'h42;
                    16'h2B18: data_out = 8'h43;
                    16'h2B19: data_out = 8'h44;
                    16'h2B1A: data_out = 8'h45;
                    16'h2B1B: data_out = 8'h46;
                    16'h2B1C: data_out = 8'h47;
                    16'h2B1D: data_out = 8'h48;
                    16'h2B1E: data_out = 8'h49;
                    16'h2B1F: data_out = 8'h4A;
                    16'h2B20: data_out = 8'h4B;
                    16'h2B21: data_out = 8'h4C;
                    16'h2B22: data_out = 8'h4D;
                    16'h2B23: data_out = 8'h4E;
                    16'h2B24: data_out = 8'h4F;
                    16'h2B25: data_out = 8'h50;
                    16'h2B26: data_out = 8'h51;
                    16'h2B27: data_out = 8'h52;
                    16'h2B28: data_out = 8'h53;
                    16'h2B29: data_out = 8'h54;
                    16'h2B2A: data_out = 8'h55;
                    16'h2B2B: data_out = 8'h56;
                    16'h2B2C: data_out = 8'h57;
                    16'h2B2D: data_out = 8'h58;
                    16'h2B2E: data_out = 8'h59;
                    16'h2B2F: data_out = 8'h5A;
                    16'h2B30: data_out = 8'h5B;
                    16'h2B31: data_out = 8'h5C;
                    16'h2B32: data_out = 8'h5D;
                    16'h2B33: data_out = 8'h5E;
                    16'h2B34: data_out = 8'h5F;
                    16'h2B35: data_out = 8'h60;
                    16'h2B36: data_out = 8'h61;
                    16'h2B37: data_out = 8'h62;
                    16'h2B38: data_out = 8'h63;
                    16'h2B39: data_out = 8'h64;
                    16'h2B3A: data_out = 8'h65;
                    16'h2B3B: data_out = 8'h66;
                    16'h2B3C: data_out = 8'h67;
                    16'h2B3D: data_out = 8'h68;
                    16'h2B3E: data_out = 8'h69;
                    16'h2B3F: data_out = 8'h6A;
                    16'h2B40: data_out = 8'h6B;
                    16'h2B41: data_out = 8'h6C;
                    16'h2B42: data_out = 8'h6D;
                    16'h2B43: data_out = 8'h6E;
                    16'h2B44: data_out = 8'h6F;
                    16'h2B45: data_out = 8'h70;
                    16'h2B46: data_out = 8'h71;
                    16'h2B47: data_out = 8'h72;
                    16'h2B48: data_out = 8'h73;
                    16'h2B49: data_out = 8'h74;
                    16'h2B4A: data_out = 8'h75;
                    16'h2B4B: data_out = 8'h76;
                    16'h2B4C: data_out = 8'h77;
                    16'h2B4D: data_out = 8'h78;
                    16'h2B4E: data_out = 8'h79;
                    16'h2B4F: data_out = 8'h7A;
                    16'h2B50: data_out = 8'h7B;
                    16'h2B51: data_out = 8'h7C;
                    16'h2B52: data_out = 8'h7D;
                    16'h2B53: data_out = 8'h7E;
                    16'h2B54: data_out = 8'h7F;
                    16'h2B55: data_out = 8'h80;
                    16'h2B56: data_out = 8'h81;
                    16'h2B57: data_out = 8'h82;
                    16'h2B58: data_out = 8'h83;
                    16'h2B59: data_out = 8'h84;
                    16'h2B5A: data_out = 8'h85;
                    16'h2B5B: data_out = 8'h86;
                    16'h2B5C: data_out = 8'h87;
                    16'h2B5D: data_out = 8'h88;
                    16'h2B5E: data_out = 8'h89;
                    16'h2B5F: data_out = 8'h8A;
                    16'h2B60: data_out = 8'h8B;
                    16'h2B61: data_out = 8'h8C;
                    16'h2B62: data_out = 8'h8D;
                    16'h2B63: data_out = 8'h8E;
                    16'h2B64: data_out = 8'h8F;
                    16'h2B65: data_out = 8'h90;
                    16'h2B66: data_out = 8'h91;
                    16'h2B67: data_out = 8'h92;
                    16'h2B68: data_out = 8'h93;
                    16'h2B69: data_out = 8'h94;
                    16'h2B6A: data_out = 8'h95;
                    16'h2B6B: data_out = 8'h96;
                    16'h2B6C: data_out = 8'h97;
                    16'h2B6D: data_out = 8'h98;
                    16'h2B6E: data_out = 8'h99;
                    16'h2B6F: data_out = 8'h9A;
                    16'h2B70: data_out = 8'h9B;
                    16'h2B71: data_out = 8'h9C;
                    16'h2B72: data_out = 8'h9D;
                    16'h2B73: data_out = 8'h9E;
                    16'h2B74: data_out = 8'h9F;
                    16'h2B75: data_out = 8'hA0;
                    16'h2B76: data_out = 8'hA1;
                    16'h2B77: data_out = 8'hA2;
                    16'h2B78: data_out = 8'hA3;
                    16'h2B79: data_out = 8'hA4;
                    16'h2B7A: data_out = 8'hA5;
                    16'h2B7B: data_out = 8'hA6;
                    16'h2B7C: data_out = 8'hA7;
                    16'h2B7D: data_out = 8'hA8;
                    16'h2B7E: data_out = 8'hA9;
                    16'h2B7F: data_out = 8'hAA;
                    16'h2B80: data_out = 8'h2B;
                    16'h2B81: data_out = 8'h2A;
                    16'h2B82: data_out = 8'h29;
                    16'h2B83: data_out = 8'h28;
                    16'h2B84: data_out = 8'h27;
                    16'h2B85: data_out = 8'h26;
                    16'h2B86: data_out = 8'h25;
                    16'h2B87: data_out = 8'h24;
                    16'h2B88: data_out = 8'h23;
                    16'h2B89: data_out = 8'h22;
                    16'h2B8A: data_out = 8'h21;
                    16'h2B8B: data_out = 8'h20;
                    16'h2B8C: data_out = 8'h1F;
                    16'h2B8D: data_out = 8'h1E;
                    16'h2B8E: data_out = 8'h1D;
                    16'h2B8F: data_out = 8'h1C;
                    16'h2B90: data_out = 8'h1B;
                    16'h2B91: data_out = 8'h1A;
                    16'h2B92: data_out = 8'h19;
                    16'h2B93: data_out = 8'h18;
                    16'h2B94: data_out = 8'h17;
                    16'h2B95: data_out = 8'h16;
                    16'h2B96: data_out = 8'h15;
                    16'h2B97: data_out = 8'h14;
                    16'h2B98: data_out = 8'h13;
                    16'h2B99: data_out = 8'h12;
                    16'h2B9A: data_out = 8'h11;
                    16'h2B9B: data_out = 8'h10;
                    16'h2B9C: data_out = 8'hF;
                    16'h2B9D: data_out = 8'hE;
                    16'h2B9E: data_out = 8'hD;
                    16'h2B9F: data_out = 8'hC;
                    16'h2BA0: data_out = 8'hB;
                    16'h2BA1: data_out = 8'hA;
                    16'h2BA2: data_out = 8'h9;
                    16'h2BA3: data_out = 8'h8;
                    16'h2BA4: data_out = 8'h7;
                    16'h2BA5: data_out = 8'h6;
                    16'h2BA6: data_out = 8'h5;
                    16'h2BA7: data_out = 8'h4;
                    16'h2BA8: data_out = 8'h3;
                    16'h2BA9: data_out = 8'h2;
                    16'h2BAA: data_out = 8'h1;
                    16'h2BAB: data_out = 8'h0;
                    16'h2BAC: data_out = 8'h81;
                    16'h2BAD: data_out = 8'h82;
                    16'h2BAE: data_out = 8'h83;
                    16'h2BAF: data_out = 8'h84;
                    16'h2BB0: data_out = 8'h85;
                    16'h2BB1: data_out = 8'h86;
                    16'h2BB2: data_out = 8'h87;
                    16'h2BB3: data_out = 8'h88;
                    16'h2BB4: data_out = 8'h89;
                    16'h2BB5: data_out = 8'h8A;
                    16'h2BB6: data_out = 8'h8B;
                    16'h2BB7: data_out = 8'h8C;
                    16'h2BB8: data_out = 8'h8D;
                    16'h2BB9: data_out = 8'h8E;
                    16'h2BBA: data_out = 8'h8F;
                    16'h2BBB: data_out = 8'h90;
                    16'h2BBC: data_out = 8'h91;
                    16'h2BBD: data_out = 8'h92;
                    16'h2BBE: data_out = 8'h93;
                    16'h2BBF: data_out = 8'h94;
                    16'h2BC0: data_out = 8'h95;
                    16'h2BC1: data_out = 8'h96;
                    16'h2BC2: data_out = 8'h97;
                    16'h2BC3: data_out = 8'h98;
                    16'h2BC4: data_out = 8'h99;
                    16'h2BC5: data_out = 8'h9A;
                    16'h2BC6: data_out = 8'h9B;
                    16'h2BC7: data_out = 8'h9C;
                    16'h2BC8: data_out = 8'h9D;
                    16'h2BC9: data_out = 8'h9E;
                    16'h2BCA: data_out = 8'h9F;
                    16'h2BCB: data_out = 8'hA0;
                    16'h2BCC: data_out = 8'hA1;
                    16'h2BCD: data_out = 8'hA2;
                    16'h2BCE: data_out = 8'hA3;
                    16'h2BCF: data_out = 8'hA4;
                    16'h2BD0: data_out = 8'hA5;
                    16'h2BD1: data_out = 8'hA6;
                    16'h2BD2: data_out = 8'hA7;
                    16'h2BD3: data_out = 8'hA8;
                    16'h2BD4: data_out = 8'hA9;
                    16'h2BD5: data_out = 8'hAA;
                    16'h2BD6: data_out = 8'hAB;
                    16'h2BD7: data_out = 8'hAC;
                    16'h2BD8: data_out = 8'hAD;
                    16'h2BD9: data_out = 8'hAE;
                    16'h2BDA: data_out = 8'hAF;
                    16'h2BDB: data_out = 8'hB0;
                    16'h2BDC: data_out = 8'hB1;
                    16'h2BDD: data_out = 8'hB2;
                    16'h2BDE: data_out = 8'hB3;
                    16'h2BDF: data_out = 8'hB4;
                    16'h2BE0: data_out = 8'hB5;
                    16'h2BE1: data_out = 8'hB6;
                    16'h2BE2: data_out = 8'hB7;
                    16'h2BE3: data_out = 8'hB8;
                    16'h2BE4: data_out = 8'hB9;
                    16'h2BE5: data_out = 8'hBA;
                    16'h2BE6: data_out = 8'hBB;
                    16'h2BE7: data_out = 8'hBC;
                    16'h2BE8: data_out = 8'hBD;
                    16'h2BE9: data_out = 8'hBE;
                    16'h2BEA: data_out = 8'hBF;
                    16'h2BEB: data_out = 8'hC0;
                    16'h2BEC: data_out = 8'hC1;
                    16'h2BED: data_out = 8'hC2;
                    16'h2BEE: data_out = 8'hC3;
                    16'h2BEF: data_out = 8'hC4;
                    16'h2BF0: data_out = 8'hC5;
                    16'h2BF1: data_out = 8'hC6;
                    16'h2BF2: data_out = 8'hC7;
                    16'h2BF3: data_out = 8'hC8;
                    16'h2BF4: data_out = 8'hC9;
                    16'h2BF5: data_out = 8'hCA;
                    16'h2BF6: data_out = 8'hCB;
                    16'h2BF7: data_out = 8'hCC;
                    16'h2BF8: data_out = 8'hCD;
                    16'h2BF9: data_out = 8'hCE;
                    16'h2BFA: data_out = 8'hCF;
                    16'h2BFB: data_out = 8'hD0;
                    16'h2BFC: data_out = 8'hD1;
                    16'h2BFD: data_out = 8'hD2;
                    16'h2BFE: data_out = 8'hD3;
                    16'h2BFF: data_out = 8'hD4;
                    16'h2C00: data_out = 8'h2C;
                    16'h2C01: data_out = 8'h2D;
                    16'h2C02: data_out = 8'h2E;
                    16'h2C03: data_out = 8'h2F;
                    16'h2C04: data_out = 8'h30;
                    16'h2C05: data_out = 8'h31;
                    16'h2C06: data_out = 8'h32;
                    16'h2C07: data_out = 8'h33;
                    16'h2C08: data_out = 8'h34;
                    16'h2C09: data_out = 8'h35;
                    16'h2C0A: data_out = 8'h36;
                    16'h2C0B: data_out = 8'h37;
                    16'h2C0C: data_out = 8'h38;
                    16'h2C0D: data_out = 8'h39;
                    16'h2C0E: data_out = 8'h3A;
                    16'h2C0F: data_out = 8'h3B;
                    16'h2C10: data_out = 8'h3C;
                    16'h2C11: data_out = 8'h3D;
                    16'h2C12: data_out = 8'h3E;
                    16'h2C13: data_out = 8'h3F;
                    16'h2C14: data_out = 8'h40;
                    16'h2C15: data_out = 8'h41;
                    16'h2C16: data_out = 8'h42;
                    16'h2C17: data_out = 8'h43;
                    16'h2C18: data_out = 8'h44;
                    16'h2C19: data_out = 8'h45;
                    16'h2C1A: data_out = 8'h46;
                    16'h2C1B: data_out = 8'h47;
                    16'h2C1C: data_out = 8'h48;
                    16'h2C1D: data_out = 8'h49;
                    16'h2C1E: data_out = 8'h4A;
                    16'h2C1F: data_out = 8'h4B;
                    16'h2C20: data_out = 8'h4C;
                    16'h2C21: data_out = 8'h4D;
                    16'h2C22: data_out = 8'h4E;
                    16'h2C23: data_out = 8'h4F;
                    16'h2C24: data_out = 8'h50;
                    16'h2C25: data_out = 8'h51;
                    16'h2C26: data_out = 8'h52;
                    16'h2C27: data_out = 8'h53;
                    16'h2C28: data_out = 8'h54;
                    16'h2C29: data_out = 8'h55;
                    16'h2C2A: data_out = 8'h56;
                    16'h2C2B: data_out = 8'h57;
                    16'h2C2C: data_out = 8'h58;
                    16'h2C2D: data_out = 8'h59;
                    16'h2C2E: data_out = 8'h5A;
                    16'h2C2F: data_out = 8'h5B;
                    16'h2C30: data_out = 8'h5C;
                    16'h2C31: data_out = 8'h5D;
                    16'h2C32: data_out = 8'h5E;
                    16'h2C33: data_out = 8'h5F;
                    16'h2C34: data_out = 8'h60;
                    16'h2C35: data_out = 8'h61;
                    16'h2C36: data_out = 8'h62;
                    16'h2C37: data_out = 8'h63;
                    16'h2C38: data_out = 8'h64;
                    16'h2C39: data_out = 8'h65;
                    16'h2C3A: data_out = 8'h66;
                    16'h2C3B: data_out = 8'h67;
                    16'h2C3C: data_out = 8'h68;
                    16'h2C3D: data_out = 8'h69;
                    16'h2C3E: data_out = 8'h6A;
                    16'h2C3F: data_out = 8'h6B;
                    16'h2C40: data_out = 8'h6C;
                    16'h2C41: data_out = 8'h6D;
                    16'h2C42: data_out = 8'h6E;
                    16'h2C43: data_out = 8'h6F;
                    16'h2C44: data_out = 8'h70;
                    16'h2C45: data_out = 8'h71;
                    16'h2C46: data_out = 8'h72;
                    16'h2C47: data_out = 8'h73;
                    16'h2C48: data_out = 8'h74;
                    16'h2C49: data_out = 8'h75;
                    16'h2C4A: data_out = 8'h76;
                    16'h2C4B: data_out = 8'h77;
                    16'h2C4C: data_out = 8'h78;
                    16'h2C4D: data_out = 8'h79;
                    16'h2C4E: data_out = 8'h7A;
                    16'h2C4F: data_out = 8'h7B;
                    16'h2C50: data_out = 8'h7C;
                    16'h2C51: data_out = 8'h7D;
                    16'h2C52: data_out = 8'h7E;
                    16'h2C53: data_out = 8'h7F;
                    16'h2C54: data_out = 8'h80;
                    16'h2C55: data_out = 8'h81;
                    16'h2C56: data_out = 8'h82;
                    16'h2C57: data_out = 8'h83;
                    16'h2C58: data_out = 8'h84;
                    16'h2C59: data_out = 8'h85;
                    16'h2C5A: data_out = 8'h86;
                    16'h2C5B: data_out = 8'h87;
                    16'h2C5C: data_out = 8'h88;
                    16'h2C5D: data_out = 8'h89;
                    16'h2C5E: data_out = 8'h8A;
                    16'h2C5F: data_out = 8'h8B;
                    16'h2C60: data_out = 8'h8C;
                    16'h2C61: data_out = 8'h8D;
                    16'h2C62: data_out = 8'h8E;
                    16'h2C63: data_out = 8'h8F;
                    16'h2C64: data_out = 8'h90;
                    16'h2C65: data_out = 8'h91;
                    16'h2C66: data_out = 8'h92;
                    16'h2C67: data_out = 8'h93;
                    16'h2C68: data_out = 8'h94;
                    16'h2C69: data_out = 8'h95;
                    16'h2C6A: data_out = 8'h96;
                    16'h2C6B: data_out = 8'h97;
                    16'h2C6C: data_out = 8'h98;
                    16'h2C6D: data_out = 8'h99;
                    16'h2C6E: data_out = 8'h9A;
                    16'h2C6F: data_out = 8'h9B;
                    16'h2C70: data_out = 8'h9C;
                    16'h2C71: data_out = 8'h9D;
                    16'h2C72: data_out = 8'h9E;
                    16'h2C73: data_out = 8'h9F;
                    16'h2C74: data_out = 8'hA0;
                    16'h2C75: data_out = 8'hA1;
                    16'h2C76: data_out = 8'hA2;
                    16'h2C77: data_out = 8'hA3;
                    16'h2C78: data_out = 8'hA4;
                    16'h2C79: data_out = 8'hA5;
                    16'h2C7A: data_out = 8'hA6;
                    16'h2C7B: data_out = 8'hA7;
                    16'h2C7C: data_out = 8'hA8;
                    16'h2C7D: data_out = 8'hA9;
                    16'h2C7E: data_out = 8'hAA;
                    16'h2C7F: data_out = 8'hAB;
                    16'h2C80: data_out = 8'h2C;
                    16'h2C81: data_out = 8'h2B;
                    16'h2C82: data_out = 8'h2A;
                    16'h2C83: data_out = 8'h29;
                    16'h2C84: data_out = 8'h28;
                    16'h2C85: data_out = 8'h27;
                    16'h2C86: data_out = 8'h26;
                    16'h2C87: data_out = 8'h25;
                    16'h2C88: data_out = 8'h24;
                    16'h2C89: data_out = 8'h23;
                    16'h2C8A: data_out = 8'h22;
                    16'h2C8B: data_out = 8'h21;
                    16'h2C8C: data_out = 8'h20;
                    16'h2C8D: data_out = 8'h1F;
                    16'h2C8E: data_out = 8'h1E;
                    16'h2C8F: data_out = 8'h1D;
                    16'h2C90: data_out = 8'h1C;
                    16'h2C91: data_out = 8'h1B;
                    16'h2C92: data_out = 8'h1A;
                    16'h2C93: data_out = 8'h19;
                    16'h2C94: data_out = 8'h18;
                    16'h2C95: data_out = 8'h17;
                    16'h2C96: data_out = 8'h16;
                    16'h2C97: data_out = 8'h15;
                    16'h2C98: data_out = 8'h14;
                    16'h2C99: data_out = 8'h13;
                    16'h2C9A: data_out = 8'h12;
                    16'h2C9B: data_out = 8'h11;
                    16'h2C9C: data_out = 8'h10;
                    16'h2C9D: data_out = 8'hF;
                    16'h2C9E: data_out = 8'hE;
                    16'h2C9F: data_out = 8'hD;
                    16'h2CA0: data_out = 8'hC;
                    16'h2CA1: data_out = 8'hB;
                    16'h2CA2: data_out = 8'hA;
                    16'h2CA3: data_out = 8'h9;
                    16'h2CA4: data_out = 8'h8;
                    16'h2CA5: data_out = 8'h7;
                    16'h2CA6: data_out = 8'h6;
                    16'h2CA7: data_out = 8'h5;
                    16'h2CA8: data_out = 8'h4;
                    16'h2CA9: data_out = 8'h3;
                    16'h2CAA: data_out = 8'h2;
                    16'h2CAB: data_out = 8'h1;
                    16'h2CAC: data_out = 8'h0;
                    16'h2CAD: data_out = 8'h81;
                    16'h2CAE: data_out = 8'h82;
                    16'h2CAF: data_out = 8'h83;
                    16'h2CB0: data_out = 8'h84;
                    16'h2CB1: data_out = 8'h85;
                    16'h2CB2: data_out = 8'h86;
                    16'h2CB3: data_out = 8'h87;
                    16'h2CB4: data_out = 8'h88;
                    16'h2CB5: data_out = 8'h89;
                    16'h2CB6: data_out = 8'h8A;
                    16'h2CB7: data_out = 8'h8B;
                    16'h2CB8: data_out = 8'h8C;
                    16'h2CB9: data_out = 8'h8D;
                    16'h2CBA: data_out = 8'h8E;
                    16'h2CBB: data_out = 8'h8F;
                    16'h2CBC: data_out = 8'h90;
                    16'h2CBD: data_out = 8'h91;
                    16'h2CBE: data_out = 8'h92;
                    16'h2CBF: data_out = 8'h93;
                    16'h2CC0: data_out = 8'h94;
                    16'h2CC1: data_out = 8'h95;
                    16'h2CC2: data_out = 8'h96;
                    16'h2CC3: data_out = 8'h97;
                    16'h2CC4: data_out = 8'h98;
                    16'h2CC5: data_out = 8'h99;
                    16'h2CC6: data_out = 8'h9A;
                    16'h2CC7: data_out = 8'h9B;
                    16'h2CC8: data_out = 8'h9C;
                    16'h2CC9: data_out = 8'h9D;
                    16'h2CCA: data_out = 8'h9E;
                    16'h2CCB: data_out = 8'h9F;
                    16'h2CCC: data_out = 8'hA0;
                    16'h2CCD: data_out = 8'hA1;
                    16'h2CCE: data_out = 8'hA2;
                    16'h2CCF: data_out = 8'hA3;
                    16'h2CD0: data_out = 8'hA4;
                    16'h2CD1: data_out = 8'hA5;
                    16'h2CD2: data_out = 8'hA6;
                    16'h2CD3: data_out = 8'hA7;
                    16'h2CD4: data_out = 8'hA8;
                    16'h2CD5: data_out = 8'hA9;
                    16'h2CD6: data_out = 8'hAA;
                    16'h2CD7: data_out = 8'hAB;
                    16'h2CD8: data_out = 8'hAC;
                    16'h2CD9: data_out = 8'hAD;
                    16'h2CDA: data_out = 8'hAE;
                    16'h2CDB: data_out = 8'hAF;
                    16'h2CDC: data_out = 8'hB0;
                    16'h2CDD: data_out = 8'hB1;
                    16'h2CDE: data_out = 8'hB2;
                    16'h2CDF: data_out = 8'hB3;
                    16'h2CE0: data_out = 8'hB4;
                    16'h2CE1: data_out = 8'hB5;
                    16'h2CE2: data_out = 8'hB6;
                    16'h2CE3: data_out = 8'hB7;
                    16'h2CE4: data_out = 8'hB8;
                    16'h2CE5: data_out = 8'hB9;
                    16'h2CE6: data_out = 8'hBA;
                    16'h2CE7: data_out = 8'hBB;
                    16'h2CE8: data_out = 8'hBC;
                    16'h2CE9: data_out = 8'hBD;
                    16'h2CEA: data_out = 8'hBE;
                    16'h2CEB: data_out = 8'hBF;
                    16'h2CEC: data_out = 8'hC0;
                    16'h2CED: data_out = 8'hC1;
                    16'h2CEE: data_out = 8'hC2;
                    16'h2CEF: data_out = 8'hC3;
                    16'h2CF0: data_out = 8'hC4;
                    16'h2CF1: data_out = 8'hC5;
                    16'h2CF2: data_out = 8'hC6;
                    16'h2CF3: data_out = 8'hC7;
                    16'h2CF4: data_out = 8'hC8;
                    16'h2CF5: data_out = 8'hC9;
                    16'h2CF6: data_out = 8'hCA;
                    16'h2CF7: data_out = 8'hCB;
                    16'h2CF8: data_out = 8'hCC;
                    16'h2CF9: data_out = 8'hCD;
                    16'h2CFA: data_out = 8'hCE;
                    16'h2CFB: data_out = 8'hCF;
                    16'h2CFC: data_out = 8'hD0;
                    16'h2CFD: data_out = 8'hD1;
                    16'h2CFE: data_out = 8'hD2;
                    16'h2CFF: data_out = 8'hD3;
                    16'h2D00: data_out = 8'h2D;
                    16'h2D01: data_out = 8'h2E;
                    16'h2D02: data_out = 8'h2F;
                    16'h2D03: data_out = 8'h30;
                    16'h2D04: data_out = 8'h31;
                    16'h2D05: data_out = 8'h32;
                    16'h2D06: data_out = 8'h33;
                    16'h2D07: data_out = 8'h34;
                    16'h2D08: data_out = 8'h35;
                    16'h2D09: data_out = 8'h36;
                    16'h2D0A: data_out = 8'h37;
                    16'h2D0B: data_out = 8'h38;
                    16'h2D0C: data_out = 8'h39;
                    16'h2D0D: data_out = 8'h3A;
                    16'h2D0E: data_out = 8'h3B;
                    16'h2D0F: data_out = 8'h3C;
                    16'h2D10: data_out = 8'h3D;
                    16'h2D11: data_out = 8'h3E;
                    16'h2D12: data_out = 8'h3F;
                    16'h2D13: data_out = 8'h40;
                    16'h2D14: data_out = 8'h41;
                    16'h2D15: data_out = 8'h42;
                    16'h2D16: data_out = 8'h43;
                    16'h2D17: data_out = 8'h44;
                    16'h2D18: data_out = 8'h45;
                    16'h2D19: data_out = 8'h46;
                    16'h2D1A: data_out = 8'h47;
                    16'h2D1B: data_out = 8'h48;
                    16'h2D1C: data_out = 8'h49;
                    16'h2D1D: data_out = 8'h4A;
                    16'h2D1E: data_out = 8'h4B;
                    16'h2D1F: data_out = 8'h4C;
                    16'h2D20: data_out = 8'h4D;
                    16'h2D21: data_out = 8'h4E;
                    16'h2D22: data_out = 8'h4F;
                    16'h2D23: data_out = 8'h50;
                    16'h2D24: data_out = 8'h51;
                    16'h2D25: data_out = 8'h52;
                    16'h2D26: data_out = 8'h53;
                    16'h2D27: data_out = 8'h54;
                    16'h2D28: data_out = 8'h55;
                    16'h2D29: data_out = 8'h56;
                    16'h2D2A: data_out = 8'h57;
                    16'h2D2B: data_out = 8'h58;
                    16'h2D2C: data_out = 8'h59;
                    16'h2D2D: data_out = 8'h5A;
                    16'h2D2E: data_out = 8'h5B;
                    16'h2D2F: data_out = 8'h5C;
                    16'h2D30: data_out = 8'h5D;
                    16'h2D31: data_out = 8'h5E;
                    16'h2D32: data_out = 8'h5F;
                    16'h2D33: data_out = 8'h60;
                    16'h2D34: data_out = 8'h61;
                    16'h2D35: data_out = 8'h62;
                    16'h2D36: data_out = 8'h63;
                    16'h2D37: data_out = 8'h64;
                    16'h2D38: data_out = 8'h65;
                    16'h2D39: data_out = 8'h66;
                    16'h2D3A: data_out = 8'h67;
                    16'h2D3B: data_out = 8'h68;
                    16'h2D3C: data_out = 8'h69;
                    16'h2D3D: data_out = 8'h6A;
                    16'h2D3E: data_out = 8'h6B;
                    16'h2D3F: data_out = 8'h6C;
                    16'h2D40: data_out = 8'h6D;
                    16'h2D41: data_out = 8'h6E;
                    16'h2D42: data_out = 8'h6F;
                    16'h2D43: data_out = 8'h70;
                    16'h2D44: data_out = 8'h71;
                    16'h2D45: data_out = 8'h72;
                    16'h2D46: data_out = 8'h73;
                    16'h2D47: data_out = 8'h74;
                    16'h2D48: data_out = 8'h75;
                    16'h2D49: data_out = 8'h76;
                    16'h2D4A: data_out = 8'h77;
                    16'h2D4B: data_out = 8'h78;
                    16'h2D4C: data_out = 8'h79;
                    16'h2D4D: data_out = 8'h7A;
                    16'h2D4E: data_out = 8'h7B;
                    16'h2D4F: data_out = 8'h7C;
                    16'h2D50: data_out = 8'h7D;
                    16'h2D51: data_out = 8'h7E;
                    16'h2D52: data_out = 8'h7F;
                    16'h2D53: data_out = 8'h80;
                    16'h2D54: data_out = 8'h81;
                    16'h2D55: data_out = 8'h82;
                    16'h2D56: data_out = 8'h83;
                    16'h2D57: data_out = 8'h84;
                    16'h2D58: data_out = 8'h85;
                    16'h2D59: data_out = 8'h86;
                    16'h2D5A: data_out = 8'h87;
                    16'h2D5B: data_out = 8'h88;
                    16'h2D5C: data_out = 8'h89;
                    16'h2D5D: data_out = 8'h8A;
                    16'h2D5E: data_out = 8'h8B;
                    16'h2D5F: data_out = 8'h8C;
                    16'h2D60: data_out = 8'h8D;
                    16'h2D61: data_out = 8'h8E;
                    16'h2D62: data_out = 8'h8F;
                    16'h2D63: data_out = 8'h90;
                    16'h2D64: data_out = 8'h91;
                    16'h2D65: data_out = 8'h92;
                    16'h2D66: data_out = 8'h93;
                    16'h2D67: data_out = 8'h94;
                    16'h2D68: data_out = 8'h95;
                    16'h2D69: data_out = 8'h96;
                    16'h2D6A: data_out = 8'h97;
                    16'h2D6B: data_out = 8'h98;
                    16'h2D6C: data_out = 8'h99;
                    16'h2D6D: data_out = 8'h9A;
                    16'h2D6E: data_out = 8'h9B;
                    16'h2D6F: data_out = 8'h9C;
                    16'h2D70: data_out = 8'h9D;
                    16'h2D71: data_out = 8'h9E;
                    16'h2D72: data_out = 8'h9F;
                    16'h2D73: data_out = 8'hA0;
                    16'h2D74: data_out = 8'hA1;
                    16'h2D75: data_out = 8'hA2;
                    16'h2D76: data_out = 8'hA3;
                    16'h2D77: data_out = 8'hA4;
                    16'h2D78: data_out = 8'hA5;
                    16'h2D79: data_out = 8'hA6;
                    16'h2D7A: data_out = 8'hA7;
                    16'h2D7B: data_out = 8'hA8;
                    16'h2D7C: data_out = 8'hA9;
                    16'h2D7D: data_out = 8'hAA;
                    16'h2D7E: data_out = 8'hAB;
                    16'h2D7F: data_out = 8'hAC;
                    16'h2D80: data_out = 8'h2D;
                    16'h2D81: data_out = 8'h2C;
                    16'h2D82: data_out = 8'h2B;
                    16'h2D83: data_out = 8'h2A;
                    16'h2D84: data_out = 8'h29;
                    16'h2D85: data_out = 8'h28;
                    16'h2D86: data_out = 8'h27;
                    16'h2D87: data_out = 8'h26;
                    16'h2D88: data_out = 8'h25;
                    16'h2D89: data_out = 8'h24;
                    16'h2D8A: data_out = 8'h23;
                    16'h2D8B: data_out = 8'h22;
                    16'h2D8C: data_out = 8'h21;
                    16'h2D8D: data_out = 8'h20;
                    16'h2D8E: data_out = 8'h1F;
                    16'h2D8F: data_out = 8'h1E;
                    16'h2D90: data_out = 8'h1D;
                    16'h2D91: data_out = 8'h1C;
                    16'h2D92: data_out = 8'h1B;
                    16'h2D93: data_out = 8'h1A;
                    16'h2D94: data_out = 8'h19;
                    16'h2D95: data_out = 8'h18;
                    16'h2D96: data_out = 8'h17;
                    16'h2D97: data_out = 8'h16;
                    16'h2D98: data_out = 8'h15;
                    16'h2D99: data_out = 8'h14;
                    16'h2D9A: data_out = 8'h13;
                    16'h2D9B: data_out = 8'h12;
                    16'h2D9C: data_out = 8'h11;
                    16'h2D9D: data_out = 8'h10;
                    16'h2D9E: data_out = 8'hF;
                    16'h2D9F: data_out = 8'hE;
                    16'h2DA0: data_out = 8'hD;
                    16'h2DA1: data_out = 8'hC;
                    16'h2DA2: data_out = 8'hB;
                    16'h2DA3: data_out = 8'hA;
                    16'h2DA4: data_out = 8'h9;
                    16'h2DA5: data_out = 8'h8;
                    16'h2DA6: data_out = 8'h7;
                    16'h2DA7: data_out = 8'h6;
                    16'h2DA8: data_out = 8'h5;
                    16'h2DA9: data_out = 8'h4;
                    16'h2DAA: data_out = 8'h3;
                    16'h2DAB: data_out = 8'h2;
                    16'h2DAC: data_out = 8'h1;
                    16'h2DAD: data_out = 8'h0;
                    16'h2DAE: data_out = 8'h81;
                    16'h2DAF: data_out = 8'h82;
                    16'h2DB0: data_out = 8'h83;
                    16'h2DB1: data_out = 8'h84;
                    16'h2DB2: data_out = 8'h85;
                    16'h2DB3: data_out = 8'h86;
                    16'h2DB4: data_out = 8'h87;
                    16'h2DB5: data_out = 8'h88;
                    16'h2DB6: data_out = 8'h89;
                    16'h2DB7: data_out = 8'h8A;
                    16'h2DB8: data_out = 8'h8B;
                    16'h2DB9: data_out = 8'h8C;
                    16'h2DBA: data_out = 8'h8D;
                    16'h2DBB: data_out = 8'h8E;
                    16'h2DBC: data_out = 8'h8F;
                    16'h2DBD: data_out = 8'h90;
                    16'h2DBE: data_out = 8'h91;
                    16'h2DBF: data_out = 8'h92;
                    16'h2DC0: data_out = 8'h93;
                    16'h2DC1: data_out = 8'h94;
                    16'h2DC2: data_out = 8'h95;
                    16'h2DC3: data_out = 8'h96;
                    16'h2DC4: data_out = 8'h97;
                    16'h2DC5: data_out = 8'h98;
                    16'h2DC6: data_out = 8'h99;
                    16'h2DC7: data_out = 8'h9A;
                    16'h2DC8: data_out = 8'h9B;
                    16'h2DC9: data_out = 8'h9C;
                    16'h2DCA: data_out = 8'h9D;
                    16'h2DCB: data_out = 8'h9E;
                    16'h2DCC: data_out = 8'h9F;
                    16'h2DCD: data_out = 8'hA0;
                    16'h2DCE: data_out = 8'hA1;
                    16'h2DCF: data_out = 8'hA2;
                    16'h2DD0: data_out = 8'hA3;
                    16'h2DD1: data_out = 8'hA4;
                    16'h2DD2: data_out = 8'hA5;
                    16'h2DD3: data_out = 8'hA6;
                    16'h2DD4: data_out = 8'hA7;
                    16'h2DD5: data_out = 8'hA8;
                    16'h2DD6: data_out = 8'hA9;
                    16'h2DD7: data_out = 8'hAA;
                    16'h2DD8: data_out = 8'hAB;
                    16'h2DD9: data_out = 8'hAC;
                    16'h2DDA: data_out = 8'hAD;
                    16'h2DDB: data_out = 8'hAE;
                    16'h2DDC: data_out = 8'hAF;
                    16'h2DDD: data_out = 8'hB0;
                    16'h2DDE: data_out = 8'hB1;
                    16'h2DDF: data_out = 8'hB2;
                    16'h2DE0: data_out = 8'hB3;
                    16'h2DE1: data_out = 8'hB4;
                    16'h2DE2: data_out = 8'hB5;
                    16'h2DE3: data_out = 8'hB6;
                    16'h2DE4: data_out = 8'hB7;
                    16'h2DE5: data_out = 8'hB8;
                    16'h2DE6: data_out = 8'hB9;
                    16'h2DE7: data_out = 8'hBA;
                    16'h2DE8: data_out = 8'hBB;
                    16'h2DE9: data_out = 8'hBC;
                    16'h2DEA: data_out = 8'hBD;
                    16'h2DEB: data_out = 8'hBE;
                    16'h2DEC: data_out = 8'hBF;
                    16'h2DED: data_out = 8'hC0;
                    16'h2DEE: data_out = 8'hC1;
                    16'h2DEF: data_out = 8'hC2;
                    16'h2DF0: data_out = 8'hC3;
                    16'h2DF1: data_out = 8'hC4;
                    16'h2DF2: data_out = 8'hC5;
                    16'h2DF3: data_out = 8'hC6;
                    16'h2DF4: data_out = 8'hC7;
                    16'h2DF5: data_out = 8'hC8;
                    16'h2DF6: data_out = 8'hC9;
                    16'h2DF7: data_out = 8'hCA;
                    16'h2DF8: data_out = 8'hCB;
                    16'h2DF9: data_out = 8'hCC;
                    16'h2DFA: data_out = 8'hCD;
                    16'h2DFB: data_out = 8'hCE;
                    16'h2DFC: data_out = 8'hCF;
                    16'h2DFD: data_out = 8'hD0;
                    16'h2DFE: data_out = 8'hD1;
                    16'h2DFF: data_out = 8'hD2;
                    16'h2E00: data_out = 8'h2E;
                    16'h2E01: data_out = 8'h2F;
                    16'h2E02: data_out = 8'h30;
                    16'h2E03: data_out = 8'h31;
                    16'h2E04: data_out = 8'h32;
                    16'h2E05: data_out = 8'h33;
                    16'h2E06: data_out = 8'h34;
                    16'h2E07: data_out = 8'h35;
                    16'h2E08: data_out = 8'h36;
                    16'h2E09: data_out = 8'h37;
                    16'h2E0A: data_out = 8'h38;
                    16'h2E0B: data_out = 8'h39;
                    16'h2E0C: data_out = 8'h3A;
                    16'h2E0D: data_out = 8'h3B;
                    16'h2E0E: data_out = 8'h3C;
                    16'h2E0F: data_out = 8'h3D;
                    16'h2E10: data_out = 8'h3E;
                    16'h2E11: data_out = 8'h3F;
                    16'h2E12: data_out = 8'h40;
                    16'h2E13: data_out = 8'h41;
                    16'h2E14: data_out = 8'h42;
                    16'h2E15: data_out = 8'h43;
                    16'h2E16: data_out = 8'h44;
                    16'h2E17: data_out = 8'h45;
                    16'h2E18: data_out = 8'h46;
                    16'h2E19: data_out = 8'h47;
                    16'h2E1A: data_out = 8'h48;
                    16'h2E1B: data_out = 8'h49;
                    16'h2E1C: data_out = 8'h4A;
                    16'h2E1D: data_out = 8'h4B;
                    16'h2E1E: data_out = 8'h4C;
                    16'h2E1F: data_out = 8'h4D;
                    16'h2E20: data_out = 8'h4E;
                    16'h2E21: data_out = 8'h4F;
                    16'h2E22: data_out = 8'h50;
                    16'h2E23: data_out = 8'h51;
                    16'h2E24: data_out = 8'h52;
                    16'h2E25: data_out = 8'h53;
                    16'h2E26: data_out = 8'h54;
                    16'h2E27: data_out = 8'h55;
                    16'h2E28: data_out = 8'h56;
                    16'h2E29: data_out = 8'h57;
                    16'h2E2A: data_out = 8'h58;
                    16'h2E2B: data_out = 8'h59;
                    16'h2E2C: data_out = 8'h5A;
                    16'h2E2D: data_out = 8'h5B;
                    16'h2E2E: data_out = 8'h5C;
                    16'h2E2F: data_out = 8'h5D;
                    16'h2E30: data_out = 8'h5E;
                    16'h2E31: data_out = 8'h5F;
                    16'h2E32: data_out = 8'h60;
                    16'h2E33: data_out = 8'h61;
                    16'h2E34: data_out = 8'h62;
                    16'h2E35: data_out = 8'h63;
                    16'h2E36: data_out = 8'h64;
                    16'h2E37: data_out = 8'h65;
                    16'h2E38: data_out = 8'h66;
                    16'h2E39: data_out = 8'h67;
                    16'h2E3A: data_out = 8'h68;
                    16'h2E3B: data_out = 8'h69;
                    16'h2E3C: data_out = 8'h6A;
                    16'h2E3D: data_out = 8'h6B;
                    16'h2E3E: data_out = 8'h6C;
                    16'h2E3F: data_out = 8'h6D;
                    16'h2E40: data_out = 8'h6E;
                    16'h2E41: data_out = 8'h6F;
                    16'h2E42: data_out = 8'h70;
                    16'h2E43: data_out = 8'h71;
                    16'h2E44: data_out = 8'h72;
                    16'h2E45: data_out = 8'h73;
                    16'h2E46: data_out = 8'h74;
                    16'h2E47: data_out = 8'h75;
                    16'h2E48: data_out = 8'h76;
                    16'h2E49: data_out = 8'h77;
                    16'h2E4A: data_out = 8'h78;
                    16'h2E4B: data_out = 8'h79;
                    16'h2E4C: data_out = 8'h7A;
                    16'h2E4D: data_out = 8'h7B;
                    16'h2E4E: data_out = 8'h7C;
                    16'h2E4F: data_out = 8'h7D;
                    16'h2E50: data_out = 8'h7E;
                    16'h2E51: data_out = 8'h7F;
                    16'h2E52: data_out = 8'h80;
                    16'h2E53: data_out = 8'h81;
                    16'h2E54: data_out = 8'h82;
                    16'h2E55: data_out = 8'h83;
                    16'h2E56: data_out = 8'h84;
                    16'h2E57: data_out = 8'h85;
                    16'h2E58: data_out = 8'h86;
                    16'h2E59: data_out = 8'h87;
                    16'h2E5A: data_out = 8'h88;
                    16'h2E5B: data_out = 8'h89;
                    16'h2E5C: data_out = 8'h8A;
                    16'h2E5D: data_out = 8'h8B;
                    16'h2E5E: data_out = 8'h8C;
                    16'h2E5F: data_out = 8'h8D;
                    16'h2E60: data_out = 8'h8E;
                    16'h2E61: data_out = 8'h8F;
                    16'h2E62: data_out = 8'h90;
                    16'h2E63: data_out = 8'h91;
                    16'h2E64: data_out = 8'h92;
                    16'h2E65: data_out = 8'h93;
                    16'h2E66: data_out = 8'h94;
                    16'h2E67: data_out = 8'h95;
                    16'h2E68: data_out = 8'h96;
                    16'h2E69: data_out = 8'h97;
                    16'h2E6A: data_out = 8'h98;
                    16'h2E6B: data_out = 8'h99;
                    16'h2E6C: data_out = 8'h9A;
                    16'h2E6D: data_out = 8'h9B;
                    16'h2E6E: data_out = 8'h9C;
                    16'h2E6F: data_out = 8'h9D;
                    16'h2E70: data_out = 8'h9E;
                    16'h2E71: data_out = 8'h9F;
                    16'h2E72: data_out = 8'hA0;
                    16'h2E73: data_out = 8'hA1;
                    16'h2E74: data_out = 8'hA2;
                    16'h2E75: data_out = 8'hA3;
                    16'h2E76: data_out = 8'hA4;
                    16'h2E77: data_out = 8'hA5;
                    16'h2E78: data_out = 8'hA6;
                    16'h2E79: data_out = 8'hA7;
                    16'h2E7A: data_out = 8'hA8;
                    16'h2E7B: data_out = 8'hA9;
                    16'h2E7C: data_out = 8'hAA;
                    16'h2E7D: data_out = 8'hAB;
                    16'h2E7E: data_out = 8'hAC;
                    16'h2E7F: data_out = 8'hAD;
                    16'h2E80: data_out = 8'h2E;
                    16'h2E81: data_out = 8'h2D;
                    16'h2E82: data_out = 8'h2C;
                    16'h2E83: data_out = 8'h2B;
                    16'h2E84: data_out = 8'h2A;
                    16'h2E85: data_out = 8'h29;
                    16'h2E86: data_out = 8'h28;
                    16'h2E87: data_out = 8'h27;
                    16'h2E88: data_out = 8'h26;
                    16'h2E89: data_out = 8'h25;
                    16'h2E8A: data_out = 8'h24;
                    16'h2E8B: data_out = 8'h23;
                    16'h2E8C: data_out = 8'h22;
                    16'h2E8D: data_out = 8'h21;
                    16'h2E8E: data_out = 8'h20;
                    16'h2E8F: data_out = 8'h1F;
                    16'h2E90: data_out = 8'h1E;
                    16'h2E91: data_out = 8'h1D;
                    16'h2E92: data_out = 8'h1C;
                    16'h2E93: data_out = 8'h1B;
                    16'h2E94: data_out = 8'h1A;
                    16'h2E95: data_out = 8'h19;
                    16'h2E96: data_out = 8'h18;
                    16'h2E97: data_out = 8'h17;
                    16'h2E98: data_out = 8'h16;
                    16'h2E99: data_out = 8'h15;
                    16'h2E9A: data_out = 8'h14;
                    16'h2E9B: data_out = 8'h13;
                    16'h2E9C: data_out = 8'h12;
                    16'h2E9D: data_out = 8'h11;
                    16'h2E9E: data_out = 8'h10;
                    16'h2E9F: data_out = 8'hF;
                    16'h2EA0: data_out = 8'hE;
                    16'h2EA1: data_out = 8'hD;
                    16'h2EA2: data_out = 8'hC;
                    16'h2EA3: data_out = 8'hB;
                    16'h2EA4: data_out = 8'hA;
                    16'h2EA5: data_out = 8'h9;
                    16'h2EA6: data_out = 8'h8;
                    16'h2EA7: data_out = 8'h7;
                    16'h2EA8: data_out = 8'h6;
                    16'h2EA9: data_out = 8'h5;
                    16'h2EAA: data_out = 8'h4;
                    16'h2EAB: data_out = 8'h3;
                    16'h2EAC: data_out = 8'h2;
                    16'h2EAD: data_out = 8'h1;
                    16'h2EAE: data_out = 8'h0;
                    16'h2EAF: data_out = 8'h81;
                    16'h2EB0: data_out = 8'h82;
                    16'h2EB1: data_out = 8'h83;
                    16'h2EB2: data_out = 8'h84;
                    16'h2EB3: data_out = 8'h85;
                    16'h2EB4: data_out = 8'h86;
                    16'h2EB5: data_out = 8'h87;
                    16'h2EB6: data_out = 8'h88;
                    16'h2EB7: data_out = 8'h89;
                    16'h2EB8: data_out = 8'h8A;
                    16'h2EB9: data_out = 8'h8B;
                    16'h2EBA: data_out = 8'h8C;
                    16'h2EBB: data_out = 8'h8D;
                    16'h2EBC: data_out = 8'h8E;
                    16'h2EBD: data_out = 8'h8F;
                    16'h2EBE: data_out = 8'h90;
                    16'h2EBF: data_out = 8'h91;
                    16'h2EC0: data_out = 8'h92;
                    16'h2EC1: data_out = 8'h93;
                    16'h2EC2: data_out = 8'h94;
                    16'h2EC3: data_out = 8'h95;
                    16'h2EC4: data_out = 8'h96;
                    16'h2EC5: data_out = 8'h97;
                    16'h2EC6: data_out = 8'h98;
                    16'h2EC7: data_out = 8'h99;
                    16'h2EC8: data_out = 8'h9A;
                    16'h2EC9: data_out = 8'h9B;
                    16'h2ECA: data_out = 8'h9C;
                    16'h2ECB: data_out = 8'h9D;
                    16'h2ECC: data_out = 8'h9E;
                    16'h2ECD: data_out = 8'h9F;
                    16'h2ECE: data_out = 8'hA0;
                    16'h2ECF: data_out = 8'hA1;
                    16'h2ED0: data_out = 8'hA2;
                    16'h2ED1: data_out = 8'hA3;
                    16'h2ED2: data_out = 8'hA4;
                    16'h2ED3: data_out = 8'hA5;
                    16'h2ED4: data_out = 8'hA6;
                    16'h2ED5: data_out = 8'hA7;
                    16'h2ED6: data_out = 8'hA8;
                    16'h2ED7: data_out = 8'hA9;
                    16'h2ED8: data_out = 8'hAA;
                    16'h2ED9: data_out = 8'hAB;
                    16'h2EDA: data_out = 8'hAC;
                    16'h2EDB: data_out = 8'hAD;
                    16'h2EDC: data_out = 8'hAE;
                    16'h2EDD: data_out = 8'hAF;
                    16'h2EDE: data_out = 8'hB0;
                    16'h2EDF: data_out = 8'hB1;
                    16'h2EE0: data_out = 8'hB2;
                    16'h2EE1: data_out = 8'hB3;
                    16'h2EE2: data_out = 8'hB4;
                    16'h2EE3: data_out = 8'hB5;
                    16'h2EE4: data_out = 8'hB6;
                    16'h2EE5: data_out = 8'hB7;
                    16'h2EE6: data_out = 8'hB8;
                    16'h2EE7: data_out = 8'hB9;
                    16'h2EE8: data_out = 8'hBA;
                    16'h2EE9: data_out = 8'hBB;
                    16'h2EEA: data_out = 8'hBC;
                    16'h2EEB: data_out = 8'hBD;
                    16'h2EEC: data_out = 8'hBE;
                    16'h2EED: data_out = 8'hBF;
                    16'h2EEE: data_out = 8'hC0;
                    16'h2EEF: data_out = 8'hC1;
                    16'h2EF0: data_out = 8'hC2;
                    16'h2EF1: data_out = 8'hC3;
                    16'h2EF2: data_out = 8'hC4;
                    16'h2EF3: data_out = 8'hC5;
                    16'h2EF4: data_out = 8'hC6;
                    16'h2EF5: data_out = 8'hC7;
                    16'h2EF6: data_out = 8'hC8;
                    16'h2EF7: data_out = 8'hC9;
                    16'h2EF8: data_out = 8'hCA;
                    16'h2EF9: data_out = 8'hCB;
                    16'h2EFA: data_out = 8'hCC;
                    16'h2EFB: data_out = 8'hCD;
                    16'h2EFC: data_out = 8'hCE;
                    16'h2EFD: data_out = 8'hCF;
                    16'h2EFE: data_out = 8'hD0;
                    16'h2EFF: data_out = 8'hD1;
                    16'h2F00: data_out = 8'h2F;
                    16'h2F01: data_out = 8'h30;
                    16'h2F02: data_out = 8'h31;
                    16'h2F03: data_out = 8'h32;
                    16'h2F04: data_out = 8'h33;
                    16'h2F05: data_out = 8'h34;
                    16'h2F06: data_out = 8'h35;
                    16'h2F07: data_out = 8'h36;
                    16'h2F08: data_out = 8'h37;
                    16'h2F09: data_out = 8'h38;
                    16'h2F0A: data_out = 8'h39;
                    16'h2F0B: data_out = 8'h3A;
                    16'h2F0C: data_out = 8'h3B;
                    16'h2F0D: data_out = 8'h3C;
                    16'h2F0E: data_out = 8'h3D;
                    16'h2F0F: data_out = 8'h3E;
                    16'h2F10: data_out = 8'h3F;
                    16'h2F11: data_out = 8'h40;
                    16'h2F12: data_out = 8'h41;
                    16'h2F13: data_out = 8'h42;
                    16'h2F14: data_out = 8'h43;
                    16'h2F15: data_out = 8'h44;
                    16'h2F16: data_out = 8'h45;
                    16'h2F17: data_out = 8'h46;
                    16'h2F18: data_out = 8'h47;
                    16'h2F19: data_out = 8'h48;
                    16'h2F1A: data_out = 8'h49;
                    16'h2F1B: data_out = 8'h4A;
                    16'h2F1C: data_out = 8'h4B;
                    16'h2F1D: data_out = 8'h4C;
                    16'h2F1E: data_out = 8'h4D;
                    16'h2F1F: data_out = 8'h4E;
                    16'h2F20: data_out = 8'h4F;
                    16'h2F21: data_out = 8'h50;
                    16'h2F22: data_out = 8'h51;
                    16'h2F23: data_out = 8'h52;
                    16'h2F24: data_out = 8'h53;
                    16'h2F25: data_out = 8'h54;
                    16'h2F26: data_out = 8'h55;
                    16'h2F27: data_out = 8'h56;
                    16'h2F28: data_out = 8'h57;
                    16'h2F29: data_out = 8'h58;
                    16'h2F2A: data_out = 8'h59;
                    16'h2F2B: data_out = 8'h5A;
                    16'h2F2C: data_out = 8'h5B;
                    16'h2F2D: data_out = 8'h5C;
                    16'h2F2E: data_out = 8'h5D;
                    16'h2F2F: data_out = 8'h5E;
                    16'h2F30: data_out = 8'h5F;
                    16'h2F31: data_out = 8'h60;
                    16'h2F32: data_out = 8'h61;
                    16'h2F33: data_out = 8'h62;
                    16'h2F34: data_out = 8'h63;
                    16'h2F35: data_out = 8'h64;
                    16'h2F36: data_out = 8'h65;
                    16'h2F37: data_out = 8'h66;
                    16'h2F38: data_out = 8'h67;
                    16'h2F39: data_out = 8'h68;
                    16'h2F3A: data_out = 8'h69;
                    16'h2F3B: data_out = 8'h6A;
                    16'h2F3C: data_out = 8'h6B;
                    16'h2F3D: data_out = 8'h6C;
                    16'h2F3E: data_out = 8'h6D;
                    16'h2F3F: data_out = 8'h6E;
                    16'h2F40: data_out = 8'h6F;
                    16'h2F41: data_out = 8'h70;
                    16'h2F42: data_out = 8'h71;
                    16'h2F43: data_out = 8'h72;
                    16'h2F44: data_out = 8'h73;
                    16'h2F45: data_out = 8'h74;
                    16'h2F46: data_out = 8'h75;
                    16'h2F47: data_out = 8'h76;
                    16'h2F48: data_out = 8'h77;
                    16'h2F49: data_out = 8'h78;
                    16'h2F4A: data_out = 8'h79;
                    16'h2F4B: data_out = 8'h7A;
                    16'h2F4C: data_out = 8'h7B;
                    16'h2F4D: data_out = 8'h7C;
                    16'h2F4E: data_out = 8'h7D;
                    16'h2F4F: data_out = 8'h7E;
                    16'h2F50: data_out = 8'h7F;
                    16'h2F51: data_out = 8'h80;
                    16'h2F52: data_out = 8'h81;
                    16'h2F53: data_out = 8'h82;
                    16'h2F54: data_out = 8'h83;
                    16'h2F55: data_out = 8'h84;
                    16'h2F56: data_out = 8'h85;
                    16'h2F57: data_out = 8'h86;
                    16'h2F58: data_out = 8'h87;
                    16'h2F59: data_out = 8'h88;
                    16'h2F5A: data_out = 8'h89;
                    16'h2F5B: data_out = 8'h8A;
                    16'h2F5C: data_out = 8'h8B;
                    16'h2F5D: data_out = 8'h8C;
                    16'h2F5E: data_out = 8'h8D;
                    16'h2F5F: data_out = 8'h8E;
                    16'h2F60: data_out = 8'h8F;
                    16'h2F61: data_out = 8'h90;
                    16'h2F62: data_out = 8'h91;
                    16'h2F63: data_out = 8'h92;
                    16'h2F64: data_out = 8'h93;
                    16'h2F65: data_out = 8'h94;
                    16'h2F66: data_out = 8'h95;
                    16'h2F67: data_out = 8'h96;
                    16'h2F68: data_out = 8'h97;
                    16'h2F69: data_out = 8'h98;
                    16'h2F6A: data_out = 8'h99;
                    16'h2F6B: data_out = 8'h9A;
                    16'h2F6C: data_out = 8'h9B;
                    16'h2F6D: data_out = 8'h9C;
                    16'h2F6E: data_out = 8'h9D;
                    16'h2F6F: data_out = 8'h9E;
                    16'h2F70: data_out = 8'h9F;
                    16'h2F71: data_out = 8'hA0;
                    16'h2F72: data_out = 8'hA1;
                    16'h2F73: data_out = 8'hA2;
                    16'h2F74: data_out = 8'hA3;
                    16'h2F75: data_out = 8'hA4;
                    16'h2F76: data_out = 8'hA5;
                    16'h2F77: data_out = 8'hA6;
                    16'h2F78: data_out = 8'hA7;
                    16'h2F79: data_out = 8'hA8;
                    16'h2F7A: data_out = 8'hA9;
                    16'h2F7B: data_out = 8'hAA;
                    16'h2F7C: data_out = 8'hAB;
                    16'h2F7D: data_out = 8'hAC;
                    16'h2F7E: data_out = 8'hAD;
                    16'h2F7F: data_out = 8'hAE;
                    16'h2F80: data_out = 8'h2F;
                    16'h2F81: data_out = 8'h2E;
                    16'h2F82: data_out = 8'h2D;
                    16'h2F83: data_out = 8'h2C;
                    16'h2F84: data_out = 8'h2B;
                    16'h2F85: data_out = 8'h2A;
                    16'h2F86: data_out = 8'h29;
                    16'h2F87: data_out = 8'h28;
                    16'h2F88: data_out = 8'h27;
                    16'h2F89: data_out = 8'h26;
                    16'h2F8A: data_out = 8'h25;
                    16'h2F8B: data_out = 8'h24;
                    16'h2F8C: data_out = 8'h23;
                    16'h2F8D: data_out = 8'h22;
                    16'h2F8E: data_out = 8'h21;
                    16'h2F8F: data_out = 8'h20;
                    16'h2F90: data_out = 8'h1F;
                    16'h2F91: data_out = 8'h1E;
                    16'h2F92: data_out = 8'h1D;
                    16'h2F93: data_out = 8'h1C;
                    16'h2F94: data_out = 8'h1B;
                    16'h2F95: data_out = 8'h1A;
                    16'h2F96: data_out = 8'h19;
                    16'h2F97: data_out = 8'h18;
                    16'h2F98: data_out = 8'h17;
                    16'h2F99: data_out = 8'h16;
                    16'h2F9A: data_out = 8'h15;
                    16'h2F9B: data_out = 8'h14;
                    16'h2F9C: data_out = 8'h13;
                    16'h2F9D: data_out = 8'h12;
                    16'h2F9E: data_out = 8'h11;
                    16'h2F9F: data_out = 8'h10;
                    16'h2FA0: data_out = 8'hF;
                    16'h2FA1: data_out = 8'hE;
                    16'h2FA2: data_out = 8'hD;
                    16'h2FA3: data_out = 8'hC;
                    16'h2FA4: data_out = 8'hB;
                    16'h2FA5: data_out = 8'hA;
                    16'h2FA6: data_out = 8'h9;
                    16'h2FA7: data_out = 8'h8;
                    16'h2FA8: data_out = 8'h7;
                    16'h2FA9: data_out = 8'h6;
                    16'h2FAA: data_out = 8'h5;
                    16'h2FAB: data_out = 8'h4;
                    16'h2FAC: data_out = 8'h3;
                    16'h2FAD: data_out = 8'h2;
                    16'h2FAE: data_out = 8'h1;
                    16'h2FAF: data_out = 8'h0;
                    16'h2FB0: data_out = 8'h81;
                    16'h2FB1: data_out = 8'h82;
                    16'h2FB2: data_out = 8'h83;
                    16'h2FB3: data_out = 8'h84;
                    16'h2FB4: data_out = 8'h85;
                    16'h2FB5: data_out = 8'h86;
                    16'h2FB6: data_out = 8'h87;
                    16'h2FB7: data_out = 8'h88;
                    16'h2FB8: data_out = 8'h89;
                    16'h2FB9: data_out = 8'h8A;
                    16'h2FBA: data_out = 8'h8B;
                    16'h2FBB: data_out = 8'h8C;
                    16'h2FBC: data_out = 8'h8D;
                    16'h2FBD: data_out = 8'h8E;
                    16'h2FBE: data_out = 8'h8F;
                    16'h2FBF: data_out = 8'h90;
                    16'h2FC0: data_out = 8'h91;
                    16'h2FC1: data_out = 8'h92;
                    16'h2FC2: data_out = 8'h93;
                    16'h2FC3: data_out = 8'h94;
                    16'h2FC4: data_out = 8'h95;
                    16'h2FC5: data_out = 8'h96;
                    16'h2FC6: data_out = 8'h97;
                    16'h2FC7: data_out = 8'h98;
                    16'h2FC8: data_out = 8'h99;
                    16'h2FC9: data_out = 8'h9A;
                    16'h2FCA: data_out = 8'h9B;
                    16'h2FCB: data_out = 8'h9C;
                    16'h2FCC: data_out = 8'h9D;
                    16'h2FCD: data_out = 8'h9E;
                    16'h2FCE: data_out = 8'h9F;
                    16'h2FCF: data_out = 8'hA0;
                    16'h2FD0: data_out = 8'hA1;
                    16'h2FD1: data_out = 8'hA2;
                    16'h2FD2: data_out = 8'hA3;
                    16'h2FD3: data_out = 8'hA4;
                    16'h2FD4: data_out = 8'hA5;
                    16'h2FD5: data_out = 8'hA6;
                    16'h2FD6: data_out = 8'hA7;
                    16'h2FD7: data_out = 8'hA8;
                    16'h2FD8: data_out = 8'hA9;
                    16'h2FD9: data_out = 8'hAA;
                    16'h2FDA: data_out = 8'hAB;
                    16'h2FDB: data_out = 8'hAC;
                    16'h2FDC: data_out = 8'hAD;
                    16'h2FDD: data_out = 8'hAE;
                    16'h2FDE: data_out = 8'hAF;
                    16'h2FDF: data_out = 8'hB0;
                    16'h2FE0: data_out = 8'hB1;
                    16'h2FE1: data_out = 8'hB2;
                    16'h2FE2: data_out = 8'hB3;
                    16'h2FE3: data_out = 8'hB4;
                    16'h2FE4: data_out = 8'hB5;
                    16'h2FE5: data_out = 8'hB6;
                    16'h2FE6: data_out = 8'hB7;
                    16'h2FE7: data_out = 8'hB8;
                    16'h2FE8: data_out = 8'hB9;
                    16'h2FE9: data_out = 8'hBA;
                    16'h2FEA: data_out = 8'hBB;
                    16'h2FEB: data_out = 8'hBC;
                    16'h2FEC: data_out = 8'hBD;
                    16'h2FED: data_out = 8'hBE;
                    16'h2FEE: data_out = 8'hBF;
                    16'h2FEF: data_out = 8'hC0;
                    16'h2FF0: data_out = 8'hC1;
                    16'h2FF1: data_out = 8'hC2;
                    16'h2FF2: data_out = 8'hC3;
                    16'h2FF3: data_out = 8'hC4;
                    16'h2FF4: data_out = 8'hC5;
                    16'h2FF5: data_out = 8'hC6;
                    16'h2FF6: data_out = 8'hC7;
                    16'h2FF7: data_out = 8'hC8;
                    16'h2FF8: data_out = 8'hC9;
                    16'h2FF9: data_out = 8'hCA;
                    16'h2FFA: data_out = 8'hCB;
                    16'h2FFB: data_out = 8'hCC;
                    16'h2FFC: data_out = 8'hCD;
                    16'h2FFD: data_out = 8'hCE;
                    16'h2FFE: data_out = 8'hCF;
                    16'h2FFF: data_out = 8'hD0;
                    16'h3000: data_out = 8'h30;
                    16'h3001: data_out = 8'h31;
                    16'h3002: data_out = 8'h32;
                    16'h3003: data_out = 8'h33;
                    16'h3004: data_out = 8'h34;
                    16'h3005: data_out = 8'h35;
                    16'h3006: data_out = 8'h36;
                    16'h3007: data_out = 8'h37;
                    16'h3008: data_out = 8'h38;
                    16'h3009: data_out = 8'h39;
                    16'h300A: data_out = 8'h3A;
                    16'h300B: data_out = 8'h3B;
                    16'h300C: data_out = 8'h3C;
                    16'h300D: data_out = 8'h3D;
                    16'h300E: data_out = 8'h3E;
                    16'h300F: data_out = 8'h3F;
                    16'h3010: data_out = 8'h40;
                    16'h3011: data_out = 8'h41;
                    16'h3012: data_out = 8'h42;
                    16'h3013: data_out = 8'h43;
                    16'h3014: data_out = 8'h44;
                    16'h3015: data_out = 8'h45;
                    16'h3016: data_out = 8'h46;
                    16'h3017: data_out = 8'h47;
                    16'h3018: data_out = 8'h48;
                    16'h3019: data_out = 8'h49;
                    16'h301A: data_out = 8'h4A;
                    16'h301B: data_out = 8'h4B;
                    16'h301C: data_out = 8'h4C;
                    16'h301D: data_out = 8'h4D;
                    16'h301E: data_out = 8'h4E;
                    16'h301F: data_out = 8'h4F;
                    16'h3020: data_out = 8'h50;
                    16'h3021: data_out = 8'h51;
                    16'h3022: data_out = 8'h52;
                    16'h3023: data_out = 8'h53;
                    16'h3024: data_out = 8'h54;
                    16'h3025: data_out = 8'h55;
                    16'h3026: data_out = 8'h56;
                    16'h3027: data_out = 8'h57;
                    16'h3028: data_out = 8'h58;
                    16'h3029: data_out = 8'h59;
                    16'h302A: data_out = 8'h5A;
                    16'h302B: data_out = 8'h5B;
                    16'h302C: data_out = 8'h5C;
                    16'h302D: data_out = 8'h5D;
                    16'h302E: data_out = 8'h5E;
                    16'h302F: data_out = 8'h5F;
                    16'h3030: data_out = 8'h60;
                    16'h3031: data_out = 8'h61;
                    16'h3032: data_out = 8'h62;
                    16'h3033: data_out = 8'h63;
                    16'h3034: data_out = 8'h64;
                    16'h3035: data_out = 8'h65;
                    16'h3036: data_out = 8'h66;
                    16'h3037: data_out = 8'h67;
                    16'h3038: data_out = 8'h68;
                    16'h3039: data_out = 8'h69;
                    16'h303A: data_out = 8'h6A;
                    16'h303B: data_out = 8'h6B;
                    16'h303C: data_out = 8'h6C;
                    16'h303D: data_out = 8'h6D;
                    16'h303E: data_out = 8'h6E;
                    16'h303F: data_out = 8'h6F;
                    16'h3040: data_out = 8'h70;
                    16'h3041: data_out = 8'h71;
                    16'h3042: data_out = 8'h72;
                    16'h3043: data_out = 8'h73;
                    16'h3044: data_out = 8'h74;
                    16'h3045: data_out = 8'h75;
                    16'h3046: data_out = 8'h76;
                    16'h3047: data_out = 8'h77;
                    16'h3048: data_out = 8'h78;
                    16'h3049: data_out = 8'h79;
                    16'h304A: data_out = 8'h7A;
                    16'h304B: data_out = 8'h7B;
                    16'h304C: data_out = 8'h7C;
                    16'h304D: data_out = 8'h7D;
                    16'h304E: data_out = 8'h7E;
                    16'h304F: data_out = 8'h7F;
                    16'h3050: data_out = 8'h80;
                    16'h3051: data_out = 8'h81;
                    16'h3052: data_out = 8'h82;
                    16'h3053: data_out = 8'h83;
                    16'h3054: data_out = 8'h84;
                    16'h3055: data_out = 8'h85;
                    16'h3056: data_out = 8'h86;
                    16'h3057: data_out = 8'h87;
                    16'h3058: data_out = 8'h88;
                    16'h3059: data_out = 8'h89;
                    16'h305A: data_out = 8'h8A;
                    16'h305B: data_out = 8'h8B;
                    16'h305C: data_out = 8'h8C;
                    16'h305D: data_out = 8'h8D;
                    16'h305E: data_out = 8'h8E;
                    16'h305F: data_out = 8'h8F;
                    16'h3060: data_out = 8'h90;
                    16'h3061: data_out = 8'h91;
                    16'h3062: data_out = 8'h92;
                    16'h3063: data_out = 8'h93;
                    16'h3064: data_out = 8'h94;
                    16'h3065: data_out = 8'h95;
                    16'h3066: data_out = 8'h96;
                    16'h3067: data_out = 8'h97;
                    16'h3068: data_out = 8'h98;
                    16'h3069: data_out = 8'h99;
                    16'h306A: data_out = 8'h9A;
                    16'h306B: data_out = 8'h9B;
                    16'h306C: data_out = 8'h9C;
                    16'h306D: data_out = 8'h9D;
                    16'h306E: data_out = 8'h9E;
                    16'h306F: data_out = 8'h9F;
                    16'h3070: data_out = 8'hA0;
                    16'h3071: data_out = 8'hA1;
                    16'h3072: data_out = 8'hA2;
                    16'h3073: data_out = 8'hA3;
                    16'h3074: data_out = 8'hA4;
                    16'h3075: data_out = 8'hA5;
                    16'h3076: data_out = 8'hA6;
                    16'h3077: data_out = 8'hA7;
                    16'h3078: data_out = 8'hA8;
                    16'h3079: data_out = 8'hA9;
                    16'h307A: data_out = 8'hAA;
                    16'h307B: data_out = 8'hAB;
                    16'h307C: data_out = 8'hAC;
                    16'h307D: data_out = 8'hAD;
                    16'h307E: data_out = 8'hAE;
                    16'h307F: data_out = 8'hAF;
                    16'h3080: data_out = 8'h30;
                    16'h3081: data_out = 8'h2F;
                    16'h3082: data_out = 8'h2E;
                    16'h3083: data_out = 8'h2D;
                    16'h3084: data_out = 8'h2C;
                    16'h3085: data_out = 8'h2B;
                    16'h3086: data_out = 8'h2A;
                    16'h3087: data_out = 8'h29;
                    16'h3088: data_out = 8'h28;
                    16'h3089: data_out = 8'h27;
                    16'h308A: data_out = 8'h26;
                    16'h308B: data_out = 8'h25;
                    16'h308C: data_out = 8'h24;
                    16'h308D: data_out = 8'h23;
                    16'h308E: data_out = 8'h22;
                    16'h308F: data_out = 8'h21;
                    16'h3090: data_out = 8'h20;
                    16'h3091: data_out = 8'h1F;
                    16'h3092: data_out = 8'h1E;
                    16'h3093: data_out = 8'h1D;
                    16'h3094: data_out = 8'h1C;
                    16'h3095: data_out = 8'h1B;
                    16'h3096: data_out = 8'h1A;
                    16'h3097: data_out = 8'h19;
                    16'h3098: data_out = 8'h18;
                    16'h3099: data_out = 8'h17;
                    16'h309A: data_out = 8'h16;
                    16'h309B: data_out = 8'h15;
                    16'h309C: data_out = 8'h14;
                    16'h309D: data_out = 8'h13;
                    16'h309E: data_out = 8'h12;
                    16'h309F: data_out = 8'h11;
                    16'h30A0: data_out = 8'h10;
                    16'h30A1: data_out = 8'hF;
                    16'h30A2: data_out = 8'hE;
                    16'h30A3: data_out = 8'hD;
                    16'h30A4: data_out = 8'hC;
                    16'h30A5: data_out = 8'hB;
                    16'h30A6: data_out = 8'hA;
                    16'h30A7: data_out = 8'h9;
                    16'h30A8: data_out = 8'h8;
                    16'h30A9: data_out = 8'h7;
                    16'h30AA: data_out = 8'h6;
                    16'h30AB: data_out = 8'h5;
                    16'h30AC: data_out = 8'h4;
                    16'h30AD: data_out = 8'h3;
                    16'h30AE: data_out = 8'h2;
                    16'h30AF: data_out = 8'h1;
                    16'h30B0: data_out = 8'h0;
                    16'h30B1: data_out = 8'h81;
                    16'h30B2: data_out = 8'h82;
                    16'h30B3: data_out = 8'h83;
                    16'h30B4: data_out = 8'h84;
                    16'h30B5: data_out = 8'h85;
                    16'h30B6: data_out = 8'h86;
                    16'h30B7: data_out = 8'h87;
                    16'h30B8: data_out = 8'h88;
                    16'h30B9: data_out = 8'h89;
                    16'h30BA: data_out = 8'h8A;
                    16'h30BB: data_out = 8'h8B;
                    16'h30BC: data_out = 8'h8C;
                    16'h30BD: data_out = 8'h8D;
                    16'h30BE: data_out = 8'h8E;
                    16'h30BF: data_out = 8'h8F;
                    16'h30C0: data_out = 8'h90;
                    16'h30C1: data_out = 8'h91;
                    16'h30C2: data_out = 8'h92;
                    16'h30C3: data_out = 8'h93;
                    16'h30C4: data_out = 8'h94;
                    16'h30C5: data_out = 8'h95;
                    16'h30C6: data_out = 8'h96;
                    16'h30C7: data_out = 8'h97;
                    16'h30C8: data_out = 8'h98;
                    16'h30C9: data_out = 8'h99;
                    16'h30CA: data_out = 8'h9A;
                    16'h30CB: data_out = 8'h9B;
                    16'h30CC: data_out = 8'h9C;
                    16'h30CD: data_out = 8'h9D;
                    16'h30CE: data_out = 8'h9E;
                    16'h30CF: data_out = 8'h9F;
                    16'h30D0: data_out = 8'hA0;
                    16'h30D1: data_out = 8'hA1;
                    16'h30D2: data_out = 8'hA2;
                    16'h30D3: data_out = 8'hA3;
                    16'h30D4: data_out = 8'hA4;
                    16'h30D5: data_out = 8'hA5;
                    16'h30D6: data_out = 8'hA6;
                    16'h30D7: data_out = 8'hA7;
                    16'h30D8: data_out = 8'hA8;
                    16'h30D9: data_out = 8'hA9;
                    16'h30DA: data_out = 8'hAA;
                    16'h30DB: data_out = 8'hAB;
                    16'h30DC: data_out = 8'hAC;
                    16'h30DD: data_out = 8'hAD;
                    16'h30DE: data_out = 8'hAE;
                    16'h30DF: data_out = 8'hAF;
                    16'h30E0: data_out = 8'hB0;
                    16'h30E1: data_out = 8'hB1;
                    16'h30E2: data_out = 8'hB2;
                    16'h30E3: data_out = 8'hB3;
                    16'h30E4: data_out = 8'hB4;
                    16'h30E5: data_out = 8'hB5;
                    16'h30E6: data_out = 8'hB6;
                    16'h30E7: data_out = 8'hB7;
                    16'h30E8: data_out = 8'hB8;
                    16'h30E9: data_out = 8'hB9;
                    16'h30EA: data_out = 8'hBA;
                    16'h30EB: data_out = 8'hBB;
                    16'h30EC: data_out = 8'hBC;
                    16'h30ED: data_out = 8'hBD;
                    16'h30EE: data_out = 8'hBE;
                    16'h30EF: data_out = 8'hBF;
                    16'h30F0: data_out = 8'hC0;
                    16'h30F1: data_out = 8'hC1;
                    16'h30F2: data_out = 8'hC2;
                    16'h30F3: data_out = 8'hC3;
                    16'h30F4: data_out = 8'hC4;
                    16'h30F5: data_out = 8'hC5;
                    16'h30F6: data_out = 8'hC6;
                    16'h30F7: data_out = 8'hC7;
                    16'h30F8: data_out = 8'hC8;
                    16'h30F9: data_out = 8'hC9;
                    16'h30FA: data_out = 8'hCA;
                    16'h30FB: data_out = 8'hCB;
                    16'h30FC: data_out = 8'hCC;
                    16'h30FD: data_out = 8'hCD;
                    16'h30FE: data_out = 8'hCE;
                    16'h30FF: data_out = 8'hCF;
                    16'h3100: data_out = 8'h31;
                    16'h3101: data_out = 8'h32;
                    16'h3102: data_out = 8'h33;
                    16'h3103: data_out = 8'h34;
                    16'h3104: data_out = 8'h35;
                    16'h3105: data_out = 8'h36;
                    16'h3106: data_out = 8'h37;
                    16'h3107: data_out = 8'h38;
                    16'h3108: data_out = 8'h39;
                    16'h3109: data_out = 8'h3A;
                    16'h310A: data_out = 8'h3B;
                    16'h310B: data_out = 8'h3C;
                    16'h310C: data_out = 8'h3D;
                    16'h310D: data_out = 8'h3E;
                    16'h310E: data_out = 8'h3F;
                    16'h310F: data_out = 8'h40;
                    16'h3110: data_out = 8'h41;
                    16'h3111: data_out = 8'h42;
                    16'h3112: data_out = 8'h43;
                    16'h3113: data_out = 8'h44;
                    16'h3114: data_out = 8'h45;
                    16'h3115: data_out = 8'h46;
                    16'h3116: data_out = 8'h47;
                    16'h3117: data_out = 8'h48;
                    16'h3118: data_out = 8'h49;
                    16'h3119: data_out = 8'h4A;
                    16'h311A: data_out = 8'h4B;
                    16'h311B: data_out = 8'h4C;
                    16'h311C: data_out = 8'h4D;
                    16'h311D: data_out = 8'h4E;
                    16'h311E: data_out = 8'h4F;
                    16'h311F: data_out = 8'h50;
                    16'h3120: data_out = 8'h51;
                    16'h3121: data_out = 8'h52;
                    16'h3122: data_out = 8'h53;
                    16'h3123: data_out = 8'h54;
                    16'h3124: data_out = 8'h55;
                    16'h3125: data_out = 8'h56;
                    16'h3126: data_out = 8'h57;
                    16'h3127: data_out = 8'h58;
                    16'h3128: data_out = 8'h59;
                    16'h3129: data_out = 8'h5A;
                    16'h312A: data_out = 8'h5B;
                    16'h312B: data_out = 8'h5C;
                    16'h312C: data_out = 8'h5D;
                    16'h312D: data_out = 8'h5E;
                    16'h312E: data_out = 8'h5F;
                    16'h312F: data_out = 8'h60;
                    16'h3130: data_out = 8'h61;
                    16'h3131: data_out = 8'h62;
                    16'h3132: data_out = 8'h63;
                    16'h3133: data_out = 8'h64;
                    16'h3134: data_out = 8'h65;
                    16'h3135: data_out = 8'h66;
                    16'h3136: data_out = 8'h67;
                    16'h3137: data_out = 8'h68;
                    16'h3138: data_out = 8'h69;
                    16'h3139: data_out = 8'h6A;
                    16'h313A: data_out = 8'h6B;
                    16'h313B: data_out = 8'h6C;
                    16'h313C: data_out = 8'h6D;
                    16'h313D: data_out = 8'h6E;
                    16'h313E: data_out = 8'h6F;
                    16'h313F: data_out = 8'h70;
                    16'h3140: data_out = 8'h71;
                    16'h3141: data_out = 8'h72;
                    16'h3142: data_out = 8'h73;
                    16'h3143: data_out = 8'h74;
                    16'h3144: data_out = 8'h75;
                    16'h3145: data_out = 8'h76;
                    16'h3146: data_out = 8'h77;
                    16'h3147: data_out = 8'h78;
                    16'h3148: data_out = 8'h79;
                    16'h3149: data_out = 8'h7A;
                    16'h314A: data_out = 8'h7B;
                    16'h314B: data_out = 8'h7C;
                    16'h314C: data_out = 8'h7D;
                    16'h314D: data_out = 8'h7E;
                    16'h314E: data_out = 8'h7F;
                    16'h314F: data_out = 8'h80;
                    16'h3150: data_out = 8'h81;
                    16'h3151: data_out = 8'h82;
                    16'h3152: data_out = 8'h83;
                    16'h3153: data_out = 8'h84;
                    16'h3154: data_out = 8'h85;
                    16'h3155: data_out = 8'h86;
                    16'h3156: data_out = 8'h87;
                    16'h3157: data_out = 8'h88;
                    16'h3158: data_out = 8'h89;
                    16'h3159: data_out = 8'h8A;
                    16'h315A: data_out = 8'h8B;
                    16'h315B: data_out = 8'h8C;
                    16'h315C: data_out = 8'h8D;
                    16'h315D: data_out = 8'h8E;
                    16'h315E: data_out = 8'h8F;
                    16'h315F: data_out = 8'h90;
                    16'h3160: data_out = 8'h91;
                    16'h3161: data_out = 8'h92;
                    16'h3162: data_out = 8'h93;
                    16'h3163: data_out = 8'h94;
                    16'h3164: data_out = 8'h95;
                    16'h3165: data_out = 8'h96;
                    16'h3166: data_out = 8'h97;
                    16'h3167: data_out = 8'h98;
                    16'h3168: data_out = 8'h99;
                    16'h3169: data_out = 8'h9A;
                    16'h316A: data_out = 8'h9B;
                    16'h316B: data_out = 8'h9C;
                    16'h316C: data_out = 8'h9D;
                    16'h316D: data_out = 8'h9E;
                    16'h316E: data_out = 8'h9F;
                    16'h316F: data_out = 8'hA0;
                    16'h3170: data_out = 8'hA1;
                    16'h3171: data_out = 8'hA2;
                    16'h3172: data_out = 8'hA3;
                    16'h3173: data_out = 8'hA4;
                    16'h3174: data_out = 8'hA5;
                    16'h3175: data_out = 8'hA6;
                    16'h3176: data_out = 8'hA7;
                    16'h3177: data_out = 8'hA8;
                    16'h3178: data_out = 8'hA9;
                    16'h3179: data_out = 8'hAA;
                    16'h317A: data_out = 8'hAB;
                    16'h317B: data_out = 8'hAC;
                    16'h317C: data_out = 8'hAD;
                    16'h317D: data_out = 8'hAE;
                    16'h317E: data_out = 8'hAF;
                    16'h317F: data_out = 8'hB0;
                    16'h3180: data_out = 8'h31;
                    16'h3181: data_out = 8'h30;
                    16'h3182: data_out = 8'h2F;
                    16'h3183: data_out = 8'h2E;
                    16'h3184: data_out = 8'h2D;
                    16'h3185: data_out = 8'h2C;
                    16'h3186: data_out = 8'h2B;
                    16'h3187: data_out = 8'h2A;
                    16'h3188: data_out = 8'h29;
                    16'h3189: data_out = 8'h28;
                    16'h318A: data_out = 8'h27;
                    16'h318B: data_out = 8'h26;
                    16'h318C: data_out = 8'h25;
                    16'h318D: data_out = 8'h24;
                    16'h318E: data_out = 8'h23;
                    16'h318F: data_out = 8'h22;
                    16'h3190: data_out = 8'h21;
                    16'h3191: data_out = 8'h20;
                    16'h3192: data_out = 8'h1F;
                    16'h3193: data_out = 8'h1E;
                    16'h3194: data_out = 8'h1D;
                    16'h3195: data_out = 8'h1C;
                    16'h3196: data_out = 8'h1B;
                    16'h3197: data_out = 8'h1A;
                    16'h3198: data_out = 8'h19;
                    16'h3199: data_out = 8'h18;
                    16'h319A: data_out = 8'h17;
                    16'h319B: data_out = 8'h16;
                    16'h319C: data_out = 8'h15;
                    16'h319D: data_out = 8'h14;
                    16'h319E: data_out = 8'h13;
                    16'h319F: data_out = 8'h12;
                    16'h31A0: data_out = 8'h11;
                    16'h31A1: data_out = 8'h10;
                    16'h31A2: data_out = 8'hF;
                    16'h31A3: data_out = 8'hE;
                    16'h31A4: data_out = 8'hD;
                    16'h31A5: data_out = 8'hC;
                    16'h31A6: data_out = 8'hB;
                    16'h31A7: data_out = 8'hA;
                    16'h31A8: data_out = 8'h9;
                    16'h31A9: data_out = 8'h8;
                    16'h31AA: data_out = 8'h7;
                    16'h31AB: data_out = 8'h6;
                    16'h31AC: data_out = 8'h5;
                    16'h31AD: data_out = 8'h4;
                    16'h31AE: data_out = 8'h3;
                    16'h31AF: data_out = 8'h2;
                    16'h31B0: data_out = 8'h1;
                    16'h31B1: data_out = 8'h0;
                    16'h31B2: data_out = 8'h81;
                    16'h31B3: data_out = 8'h82;
                    16'h31B4: data_out = 8'h83;
                    16'h31B5: data_out = 8'h84;
                    16'h31B6: data_out = 8'h85;
                    16'h31B7: data_out = 8'h86;
                    16'h31B8: data_out = 8'h87;
                    16'h31B9: data_out = 8'h88;
                    16'h31BA: data_out = 8'h89;
                    16'h31BB: data_out = 8'h8A;
                    16'h31BC: data_out = 8'h8B;
                    16'h31BD: data_out = 8'h8C;
                    16'h31BE: data_out = 8'h8D;
                    16'h31BF: data_out = 8'h8E;
                    16'h31C0: data_out = 8'h8F;
                    16'h31C1: data_out = 8'h90;
                    16'h31C2: data_out = 8'h91;
                    16'h31C3: data_out = 8'h92;
                    16'h31C4: data_out = 8'h93;
                    16'h31C5: data_out = 8'h94;
                    16'h31C6: data_out = 8'h95;
                    16'h31C7: data_out = 8'h96;
                    16'h31C8: data_out = 8'h97;
                    16'h31C9: data_out = 8'h98;
                    16'h31CA: data_out = 8'h99;
                    16'h31CB: data_out = 8'h9A;
                    16'h31CC: data_out = 8'h9B;
                    16'h31CD: data_out = 8'h9C;
                    16'h31CE: data_out = 8'h9D;
                    16'h31CF: data_out = 8'h9E;
                    16'h31D0: data_out = 8'h9F;
                    16'h31D1: data_out = 8'hA0;
                    16'h31D2: data_out = 8'hA1;
                    16'h31D3: data_out = 8'hA2;
                    16'h31D4: data_out = 8'hA3;
                    16'h31D5: data_out = 8'hA4;
                    16'h31D6: data_out = 8'hA5;
                    16'h31D7: data_out = 8'hA6;
                    16'h31D8: data_out = 8'hA7;
                    16'h31D9: data_out = 8'hA8;
                    16'h31DA: data_out = 8'hA9;
                    16'h31DB: data_out = 8'hAA;
                    16'h31DC: data_out = 8'hAB;
                    16'h31DD: data_out = 8'hAC;
                    16'h31DE: data_out = 8'hAD;
                    16'h31DF: data_out = 8'hAE;
                    16'h31E0: data_out = 8'hAF;
                    16'h31E1: data_out = 8'hB0;
                    16'h31E2: data_out = 8'hB1;
                    16'h31E3: data_out = 8'hB2;
                    16'h31E4: data_out = 8'hB3;
                    16'h31E5: data_out = 8'hB4;
                    16'h31E6: data_out = 8'hB5;
                    16'h31E7: data_out = 8'hB6;
                    16'h31E8: data_out = 8'hB7;
                    16'h31E9: data_out = 8'hB8;
                    16'h31EA: data_out = 8'hB9;
                    16'h31EB: data_out = 8'hBA;
                    16'h31EC: data_out = 8'hBB;
                    16'h31ED: data_out = 8'hBC;
                    16'h31EE: data_out = 8'hBD;
                    16'h31EF: data_out = 8'hBE;
                    16'h31F0: data_out = 8'hBF;
                    16'h31F1: data_out = 8'hC0;
                    16'h31F2: data_out = 8'hC1;
                    16'h31F3: data_out = 8'hC2;
                    16'h31F4: data_out = 8'hC3;
                    16'h31F5: data_out = 8'hC4;
                    16'h31F6: data_out = 8'hC5;
                    16'h31F7: data_out = 8'hC6;
                    16'h31F8: data_out = 8'hC7;
                    16'h31F9: data_out = 8'hC8;
                    16'h31FA: data_out = 8'hC9;
                    16'h31FB: data_out = 8'hCA;
                    16'h31FC: data_out = 8'hCB;
                    16'h31FD: data_out = 8'hCC;
                    16'h31FE: data_out = 8'hCD;
                    16'h31FF: data_out = 8'hCE;
                    16'h3200: data_out = 8'h32;
                    16'h3201: data_out = 8'h33;
                    16'h3202: data_out = 8'h34;
                    16'h3203: data_out = 8'h35;
                    16'h3204: data_out = 8'h36;
                    16'h3205: data_out = 8'h37;
                    16'h3206: data_out = 8'h38;
                    16'h3207: data_out = 8'h39;
                    16'h3208: data_out = 8'h3A;
                    16'h3209: data_out = 8'h3B;
                    16'h320A: data_out = 8'h3C;
                    16'h320B: data_out = 8'h3D;
                    16'h320C: data_out = 8'h3E;
                    16'h320D: data_out = 8'h3F;
                    16'h320E: data_out = 8'h40;
                    16'h320F: data_out = 8'h41;
                    16'h3210: data_out = 8'h42;
                    16'h3211: data_out = 8'h43;
                    16'h3212: data_out = 8'h44;
                    16'h3213: data_out = 8'h45;
                    16'h3214: data_out = 8'h46;
                    16'h3215: data_out = 8'h47;
                    16'h3216: data_out = 8'h48;
                    16'h3217: data_out = 8'h49;
                    16'h3218: data_out = 8'h4A;
                    16'h3219: data_out = 8'h4B;
                    16'h321A: data_out = 8'h4C;
                    16'h321B: data_out = 8'h4D;
                    16'h321C: data_out = 8'h4E;
                    16'h321D: data_out = 8'h4F;
                    16'h321E: data_out = 8'h50;
                    16'h321F: data_out = 8'h51;
                    16'h3220: data_out = 8'h52;
                    16'h3221: data_out = 8'h53;
                    16'h3222: data_out = 8'h54;
                    16'h3223: data_out = 8'h55;
                    16'h3224: data_out = 8'h56;
                    16'h3225: data_out = 8'h57;
                    16'h3226: data_out = 8'h58;
                    16'h3227: data_out = 8'h59;
                    16'h3228: data_out = 8'h5A;
                    16'h3229: data_out = 8'h5B;
                    16'h322A: data_out = 8'h5C;
                    16'h322B: data_out = 8'h5D;
                    16'h322C: data_out = 8'h5E;
                    16'h322D: data_out = 8'h5F;
                    16'h322E: data_out = 8'h60;
                    16'h322F: data_out = 8'h61;
                    16'h3230: data_out = 8'h62;
                    16'h3231: data_out = 8'h63;
                    16'h3232: data_out = 8'h64;
                    16'h3233: data_out = 8'h65;
                    16'h3234: data_out = 8'h66;
                    16'h3235: data_out = 8'h67;
                    16'h3236: data_out = 8'h68;
                    16'h3237: data_out = 8'h69;
                    16'h3238: data_out = 8'h6A;
                    16'h3239: data_out = 8'h6B;
                    16'h323A: data_out = 8'h6C;
                    16'h323B: data_out = 8'h6D;
                    16'h323C: data_out = 8'h6E;
                    16'h323D: data_out = 8'h6F;
                    16'h323E: data_out = 8'h70;
                    16'h323F: data_out = 8'h71;
                    16'h3240: data_out = 8'h72;
                    16'h3241: data_out = 8'h73;
                    16'h3242: data_out = 8'h74;
                    16'h3243: data_out = 8'h75;
                    16'h3244: data_out = 8'h76;
                    16'h3245: data_out = 8'h77;
                    16'h3246: data_out = 8'h78;
                    16'h3247: data_out = 8'h79;
                    16'h3248: data_out = 8'h7A;
                    16'h3249: data_out = 8'h7B;
                    16'h324A: data_out = 8'h7C;
                    16'h324B: data_out = 8'h7D;
                    16'h324C: data_out = 8'h7E;
                    16'h324D: data_out = 8'h7F;
                    16'h324E: data_out = 8'h80;
                    16'h324F: data_out = 8'h81;
                    16'h3250: data_out = 8'h82;
                    16'h3251: data_out = 8'h83;
                    16'h3252: data_out = 8'h84;
                    16'h3253: data_out = 8'h85;
                    16'h3254: data_out = 8'h86;
                    16'h3255: data_out = 8'h87;
                    16'h3256: data_out = 8'h88;
                    16'h3257: data_out = 8'h89;
                    16'h3258: data_out = 8'h8A;
                    16'h3259: data_out = 8'h8B;
                    16'h325A: data_out = 8'h8C;
                    16'h325B: data_out = 8'h8D;
                    16'h325C: data_out = 8'h8E;
                    16'h325D: data_out = 8'h8F;
                    16'h325E: data_out = 8'h90;
                    16'h325F: data_out = 8'h91;
                    16'h3260: data_out = 8'h92;
                    16'h3261: data_out = 8'h93;
                    16'h3262: data_out = 8'h94;
                    16'h3263: data_out = 8'h95;
                    16'h3264: data_out = 8'h96;
                    16'h3265: data_out = 8'h97;
                    16'h3266: data_out = 8'h98;
                    16'h3267: data_out = 8'h99;
                    16'h3268: data_out = 8'h9A;
                    16'h3269: data_out = 8'h9B;
                    16'h326A: data_out = 8'h9C;
                    16'h326B: data_out = 8'h9D;
                    16'h326C: data_out = 8'h9E;
                    16'h326D: data_out = 8'h9F;
                    16'h326E: data_out = 8'hA0;
                    16'h326F: data_out = 8'hA1;
                    16'h3270: data_out = 8'hA2;
                    16'h3271: data_out = 8'hA3;
                    16'h3272: data_out = 8'hA4;
                    16'h3273: data_out = 8'hA5;
                    16'h3274: data_out = 8'hA6;
                    16'h3275: data_out = 8'hA7;
                    16'h3276: data_out = 8'hA8;
                    16'h3277: data_out = 8'hA9;
                    16'h3278: data_out = 8'hAA;
                    16'h3279: data_out = 8'hAB;
                    16'h327A: data_out = 8'hAC;
                    16'h327B: data_out = 8'hAD;
                    16'h327C: data_out = 8'hAE;
                    16'h327D: data_out = 8'hAF;
                    16'h327E: data_out = 8'hB0;
                    16'h327F: data_out = 8'hB1;
                    16'h3280: data_out = 8'h32;
                    16'h3281: data_out = 8'h31;
                    16'h3282: data_out = 8'h30;
                    16'h3283: data_out = 8'h2F;
                    16'h3284: data_out = 8'h2E;
                    16'h3285: data_out = 8'h2D;
                    16'h3286: data_out = 8'h2C;
                    16'h3287: data_out = 8'h2B;
                    16'h3288: data_out = 8'h2A;
                    16'h3289: data_out = 8'h29;
                    16'h328A: data_out = 8'h28;
                    16'h328B: data_out = 8'h27;
                    16'h328C: data_out = 8'h26;
                    16'h328D: data_out = 8'h25;
                    16'h328E: data_out = 8'h24;
                    16'h328F: data_out = 8'h23;
                    16'h3290: data_out = 8'h22;
                    16'h3291: data_out = 8'h21;
                    16'h3292: data_out = 8'h20;
                    16'h3293: data_out = 8'h1F;
                    16'h3294: data_out = 8'h1E;
                    16'h3295: data_out = 8'h1D;
                    16'h3296: data_out = 8'h1C;
                    16'h3297: data_out = 8'h1B;
                    16'h3298: data_out = 8'h1A;
                    16'h3299: data_out = 8'h19;
                    16'h329A: data_out = 8'h18;
                    16'h329B: data_out = 8'h17;
                    16'h329C: data_out = 8'h16;
                    16'h329D: data_out = 8'h15;
                    16'h329E: data_out = 8'h14;
                    16'h329F: data_out = 8'h13;
                    16'h32A0: data_out = 8'h12;
                    16'h32A1: data_out = 8'h11;
                    16'h32A2: data_out = 8'h10;
                    16'h32A3: data_out = 8'hF;
                    16'h32A4: data_out = 8'hE;
                    16'h32A5: data_out = 8'hD;
                    16'h32A6: data_out = 8'hC;
                    16'h32A7: data_out = 8'hB;
                    16'h32A8: data_out = 8'hA;
                    16'h32A9: data_out = 8'h9;
                    16'h32AA: data_out = 8'h8;
                    16'h32AB: data_out = 8'h7;
                    16'h32AC: data_out = 8'h6;
                    16'h32AD: data_out = 8'h5;
                    16'h32AE: data_out = 8'h4;
                    16'h32AF: data_out = 8'h3;
                    16'h32B0: data_out = 8'h2;
                    16'h32B1: data_out = 8'h1;
                    16'h32B2: data_out = 8'h0;
                    16'h32B3: data_out = 8'h81;
                    16'h32B4: data_out = 8'h82;
                    16'h32B5: data_out = 8'h83;
                    16'h32B6: data_out = 8'h84;
                    16'h32B7: data_out = 8'h85;
                    16'h32B8: data_out = 8'h86;
                    16'h32B9: data_out = 8'h87;
                    16'h32BA: data_out = 8'h88;
                    16'h32BB: data_out = 8'h89;
                    16'h32BC: data_out = 8'h8A;
                    16'h32BD: data_out = 8'h8B;
                    16'h32BE: data_out = 8'h8C;
                    16'h32BF: data_out = 8'h8D;
                    16'h32C0: data_out = 8'h8E;
                    16'h32C1: data_out = 8'h8F;
                    16'h32C2: data_out = 8'h90;
                    16'h32C3: data_out = 8'h91;
                    16'h32C4: data_out = 8'h92;
                    16'h32C5: data_out = 8'h93;
                    16'h32C6: data_out = 8'h94;
                    16'h32C7: data_out = 8'h95;
                    16'h32C8: data_out = 8'h96;
                    16'h32C9: data_out = 8'h97;
                    16'h32CA: data_out = 8'h98;
                    16'h32CB: data_out = 8'h99;
                    16'h32CC: data_out = 8'h9A;
                    16'h32CD: data_out = 8'h9B;
                    16'h32CE: data_out = 8'h9C;
                    16'h32CF: data_out = 8'h9D;
                    16'h32D0: data_out = 8'h9E;
                    16'h32D1: data_out = 8'h9F;
                    16'h32D2: data_out = 8'hA0;
                    16'h32D3: data_out = 8'hA1;
                    16'h32D4: data_out = 8'hA2;
                    16'h32D5: data_out = 8'hA3;
                    16'h32D6: data_out = 8'hA4;
                    16'h32D7: data_out = 8'hA5;
                    16'h32D8: data_out = 8'hA6;
                    16'h32D9: data_out = 8'hA7;
                    16'h32DA: data_out = 8'hA8;
                    16'h32DB: data_out = 8'hA9;
                    16'h32DC: data_out = 8'hAA;
                    16'h32DD: data_out = 8'hAB;
                    16'h32DE: data_out = 8'hAC;
                    16'h32DF: data_out = 8'hAD;
                    16'h32E0: data_out = 8'hAE;
                    16'h32E1: data_out = 8'hAF;
                    16'h32E2: data_out = 8'hB0;
                    16'h32E3: data_out = 8'hB1;
                    16'h32E4: data_out = 8'hB2;
                    16'h32E5: data_out = 8'hB3;
                    16'h32E6: data_out = 8'hB4;
                    16'h32E7: data_out = 8'hB5;
                    16'h32E8: data_out = 8'hB6;
                    16'h32E9: data_out = 8'hB7;
                    16'h32EA: data_out = 8'hB8;
                    16'h32EB: data_out = 8'hB9;
                    16'h32EC: data_out = 8'hBA;
                    16'h32ED: data_out = 8'hBB;
                    16'h32EE: data_out = 8'hBC;
                    16'h32EF: data_out = 8'hBD;
                    16'h32F0: data_out = 8'hBE;
                    16'h32F1: data_out = 8'hBF;
                    16'h32F2: data_out = 8'hC0;
                    16'h32F3: data_out = 8'hC1;
                    16'h32F4: data_out = 8'hC2;
                    16'h32F5: data_out = 8'hC3;
                    16'h32F6: data_out = 8'hC4;
                    16'h32F7: data_out = 8'hC5;
                    16'h32F8: data_out = 8'hC6;
                    16'h32F9: data_out = 8'hC7;
                    16'h32FA: data_out = 8'hC8;
                    16'h32FB: data_out = 8'hC9;
                    16'h32FC: data_out = 8'hCA;
                    16'h32FD: data_out = 8'hCB;
                    16'h32FE: data_out = 8'hCC;
                    16'h32FF: data_out = 8'hCD;
                    16'h3300: data_out = 8'h33;
                    16'h3301: data_out = 8'h34;
                    16'h3302: data_out = 8'h35;
                    16'h3303: data_out = 8'h36;
                    16'h3304: data_out = 8'h37;
                    16'h3305: data_out = 8'h38;
                    16'h3306: data_out = 8'h39;
                    16'h3307: data_out = 8'h3A;
                    16'h3308: data_out = 8'h3B;
                    16'h3309: data_out = 8'h3C;
                    16'h330A: data_out = 8'h3D;
                    16'h330B: data_out = 8'h3E;
                    16'h330C: data_out = 8'h3F;
                    16'h330D: data_out = 8'h40;
                    16'h330E: data_out = 8'h41;
                    16'h330F: data_out = 8'h42;
                    16'h3310: data_out = 8'h43;
                    16'h3311: data_out = 8'h44;
                    16'h3312: data_out = 8'h45;
                    16'h3313: data_out = 8'h46;
                    16'h3314: data_out = 8'h47;
                    16'h3315: data_out = 8'h48;
                    16'h3316: data_out = 8'h49;
                    16'h3317: data_out = 8'h4A;
                    16'h3318: data_out = 8'h4B;
                    16'h3319: data_out = 8'h4C;
                    16'h331A: data_out = 8'h4D;
                    16'h331B: data_out = 8'h4E;
                    16'h331C: data_out = 8'h4F;
                    16'h331D: data_out = 8'h50;
                    16'h331E: data_out = 8'h51;
                    16'h331F: data_out = 8'h52;
                    16'h3320: data_out = 8'h53;
                    16'h3321: data_out = 8'h54;
                    16'h3322: data_out = 8'h55;
                    16'h3323: data_out = 8'h56;
                    16'h3324: data_out = 8'h57;
                    16'h3325: data_out = 8'h58;
                    16'h3326: data_out = 8'h59;
                    16'h3327: data_out = 8'h5A;
                    16'h3328: data_out = 8'h5B;
                    16'h3329: data_out = 8'h5C;
                    16'h332A: data_out = 8'h5D;
                    16'h332B: data_out = 8'h5E;
                    16'h332C: data_out = 8'h5F;
                    16'h332D: data_out = 8'h60;
                    16'h332E: data_out = 8'h61;
                    16'h332F: data_out = 8'h62;
                    16'h3330: data_out = 8'h63;
                    16'h3331: data_out = 8'h64;
                    16'h3332: data_out = 8'h65;
                    16'h3333: data_out = 8'h66;
                    16'h3334: data_out = 8'h67;
                    16'h3335: data_out = 8'h68;
                    16'h3336: data_out = 8'h69;
                    16'h3337: data_out = 8'h6A;
                    16'h3338: data_out = 8'h6B;
                    16'h3339: data_out = 8'h6C;
                    16'h333A: data_out = 8'h6D;
                    16'h333B: data_out = 8'h6E;
                    16'h333C: data_out = 8'h6F;
                    16'h333D: data_out = 8'h70;
                    16'h333E: data_out = 8'h71;
                    16'h333F: data_out = 8'h72;
                    16'h3340: data_out = 8'h73;
                    16'h3341: data_out = 8'h74;
                    16'h3342: data_out = 8'h75;
                    16'h3343: data_out = 8'h76;
                    16'h3344: data_out = 8'h77;
                    16'h3345: data_out = 8'h78;
                    16'h3346: data_out = 8'h79;
                    16'h3347: data_out = 8'h7A;
                    16'h3348: data_out = 8'h7B;
                    16'h3349: data_out = 8'h7C;
                    16'h334A: data_out = 8'h7D;
                    16'h334B: data_out = 8'h7E;
                    16'h334C: data_out = 8'h7F;
                    16'h334D: data_out = 8'h80;
                    16'h334E: data_out = 8'h81;
                    16'h334F: data_out = 8'h82;
                    16'h3350: data_out = 8'h83;
                    16'h3351: data_out = 8'h84;
                    16'h3352: data_out = 8'h85;
                    16'h3353: data_out = 8'h86;
                    16'h3354: data_out = 8'h87;
                    16'h3355: data_out = 8'h88;
                    16'h3356: data_out = 8'h89;
                    16'h3357: data_out = 8'h8A;
                    16'h3358: data_out = 8'h8B;
                    16'h3359: data_out = 8'h8C;
                    16'h335A: data_out = 8'h8D;
                    16'h335B: data_out = 8'h8E;
                    16'h335C: data_out = 8'h8F;
                    16'h335D: data_out = 8'h90;
                    16'h335E: data_out = 8'h91;
                    16'h335F: data_out = 8'h92;
                    16'h3360: data_out = 8'h93;
                    16'h3361: data_out = 8'h94;
                    16'h3362: data_out = 8'h95;
                    16'h3363: data_out = 8'h96;
                    16'h3364: data_out = 8'h97;
                    16'h3365: data_out = 8'h98;
                    16'h3366: data_out = 8'h99;
                    16'h3367: data_out = 8'h9A;
                    16'h3368: data_out = 8'h9B;
                    16'h3369: data_out = 8'h9C;
                    16'h336A: data_out = 8'h9D;
                    16'h336B: data_out = 8'h9E;
                    16'h336C: data_out = 8'h9F;
                    16'h336D: data_out = 8'hA0;
                    16'h336E: data_out = 8'hA1;
                    16'h336F: data_out = 8'hA2;
                    16'h3370: data_out = 8'hA3;
                    16'h3371: data_out = 8'hA4;
                    16'h3372: data_out = 8'hA5;
                    16'h3373: data_out = 8'hA6;
                    16'h3374: data_out = 8'hA7;
                    16'h3375: data_out = 8'hA8;
                    16'h3376: data_out = 8'hA9;
                    16'h3377: data_out = 8'hAA;
                    16'h3378: data_out = 8'hAB;
                    16'h3379: data_out = 8'hAC;
                    16'h337A: data_out = 8'hAD;
                    16'h337B: data_out = 8'hAE;
                    16'h337C: data_out = 8'hAF;
                    16'h337D: data_out = 8'hB0;
                    16'h337E: data_out = 8'hB1;
                    16'h337F: data_out = 8'hB2;
                    16'h3380: data_out = 8'h33;
                    16'h3381: data_out = 8'h32;
                    16'h3382: data_out = 8'h31;
                    16'h3383: data_out = 8'h30;
                    16'h3384: data_out = 8'h2F;
                    16'h3385: data_out = 8'h2E;
                    16'h3386: data_out = 8'h2D;
                    16'h3387: data_out = 8'h2C;
                    16'h3388: data_out = 8'h2B;
                    16'h3389: data_out = 8'h2A;
                    16'h338A: data_out = 8'h29;
                    16'h338B: data_out = 8'h28;
                    16'h338C: data_out = 8'h27;
                    16'h338D: data_out = 8'h26;
                    16'h338E: data_out = 8'h25;
                    16'h338F: data_out = 8'h24;
                    16'h3390: data_out = 8'h23;
                    16'h3391: data_out = 8'h22;
                    16'h3392: data_out = 8'h21;
                    16'h3393: data_out = 8'h20;
                    16'h3394: data_out = 8'h1F;
                    16'h3395: data_out = 8'h1E;
                    16'h3396: data_out = 8'h1D;
                    16'h3397: data_out = 8'h1C;
                    16'h3398: data_out = 8'h1B;
                    16'h3399: data_out = 8'h1A;
                    16'h339A: data_out = 8'h19;
                    16'h339B: data_out = 8'h18;
                    16'h339C: data_out = 8'h17;
                    16'h339D: data_out = 8'h16;
                    16'h339E: data_out = 8'h15;
                    16'h339F: data_out = 8'h14;
                    16'h33A0: data_out = 8'h13;
                    16'h33A1: data_out = 8'h12;
                    16'h33A2: data_out = 8'h11;
                    16'h33A3: data_out = 8'h10;
                    16'h33A4: data_out = 8'hF;
                    16'h33A5: data_out = 8'hE;
                    16'h33A6: data_out = 8'hD;
                    16'h33A7: data_out = 8'hC;
                    16'h33A8: data_out = 8'hB;
                    16'h33A9: data_out = 8'hA;
                    16'h33AA: data_out = 8'h9;
                    16'h33AB: data_out = 8'h8;
                    16'h33AC: data_out = 8'h7;
                    16'h33AD: data_out = 8'h6;
                    16'h33AE: data_out = 8'h5;
                    16'h33AF: data_out = 8'h4;
                    16'h33B0: data_out = 8'h3;
                    16'h33B1: data_out = 8'h2;
                    16'h33B2: data_out = 8'h1;
                    16'h33B3: data_out = 8'h0;
                    16'h33B4: data_out = 8'h81;
                    16'h33B5: data_out = 8'h82;
                    16'h33B6: data_out = 8'h83;
                    16'h33B7: data_out = 8'h84;
                    16'h33B8: data_out = 8'h85;
                    16'h33B9: data_out = 8'h86;
                    16'h33BA: data_out = 8'h87;
                    16'h33BB: data_out = 8'h88;
                    16'h33BC: data_out = 8'h89;
                    16'h33BD: data_out = 8'h8A;
                    16'h33BE: data_out = 8'h8B;
                    16'h33BF: data_out = 8'h8C;
                    16'h33C0: data_out = 8'h8D;
                    16'h33C1: data_out = 8'h8E;
                    16'h33C2: data_out = 8'h8F;
                    16'h33C3: data_out = 8'h90;
                    16'h33C4: data_out = 8'h91;
                    16'h33C5: data_out = 8'h92;
                    16'h33C6: data_out = 8'h93;
                    16'h33C7: data_out = 8'h94;
                    16'h33C8: data_out = 8'h95;
                    16'h33C9: data_out = 8'h96;
                    16'h33CA: data_out = 8'h97;
                    16'h33CB: data_out = 8'h98;
                    16'h33CC: data_out = 8'h99;
                    16'h33CD: data_out = 8'h9A;
                    16'h33CE: data_out = 8'h9B;
                    16'h33CF: data_out = 8'h9C;
                    16'h33D0: data_out = 8'h9D;
                    16'h33D1: data_out = 8'h9E;
                    16'h33D2: data_out = 8'h9F;
                    16'h33D3: data_out = 8'hA0;
                    16'h33D4: data_out = 8'hA1;
                    16'h33D5: data_out = 8'hA2;
                    16'h33D6: data_out = 8'hA3;
                    16'h33D7: data_out = 8'hA4;
                    16'h33D8: data_out = 8'hA5;
                    16'h33D9: data_out = 8'hA6;
                    16'h33DA: data_out = 8'hA7;
                    16'h33DB: data_out = 8'hA8;
                    16'h33DC: data_out = 8'hA9;
                    16'h33DD: data_out = 8'hAA;
                    16'h33DE: data_out = 8'hAB;
                    16'h33DF: data_out = 8'hAC;
                    16'h33E0: data_out = 8'hAD;
                    16'h33E1: data_out = 8'hAE;
                    16'h33E2: data_out = 8'hAF;
                    16'h33E3: data_out = 8'hB0;
                    16'h33E4: data_out = 8'hB1;
                    16'h33E5: data_out = 8'hB2;
                    16'h33E6: data_out = 8'hB3;
                    16'h33E7: data_out = 8'hB4;
                    16'h33E8: data_out = 8'hB5;
                    16'h33E9: data_out = 8'hB6;
                    16'h33EA: data_out = 8'hB7;
                    16'h33EB: data_out = 8'hB8;
                    16'h33EC: data_out = 8'hB9;
                    16'h33ED: data_out = 8'hBA;
                    16'h33EE: data_out = 8'hBB;
                    16'h33EF: data_out = 8'hBC;
                    16'h33F0: data_out = 8'hBD;
                    16'h33F1: data_out = 8'hBE;
                    16'h33F2: data_out = 8'hBF;
                    16'h33F3: data_out = 8'hC0;
                    16'h33F4: data_out = 8'hC1;
                    16'h33F5: data_out = 8'hC2;
                    16'h33F6: data_out = 8'hC3;
                    16'h33F7: data_out = 8'hC4;
                    16'h33F8: data_out = 8'hC5;
                    16'h33F9: data_out = 8'hC6;
                    16'h33FA: data_out = 8'hC7;
                    16'h33FB: data_out = 8'hC8;
                    16'h33FC: data_out = 8'hC9;
                    16'h33FD: data_out = 8'hCA;
                    16'h33FE: data_out = 8'hCB;
                    16'h33FF: data_out = 8'hCC;
                    16'h3400: data_out = 8'h34;
                    16'h3401: data_out = 8'h35;
                    16'h3402: data_out = 8'h36;
                    16'h3403: data_out = 8'h37;
                    16'h3404: data_out = 8'h38;
                    16'h3405: data_out = 8'h39;
                    16'h3406: data_out = 8'h3A;
                    16'h3407: data_out = 8'h3B;
                    16'h3408: data_out = 8'h3C;
                    16'h3409: data_out = 8'h3D;
                    16'h340A: data_out = 8'h3E;
                    16'h340B: data_out = 8'h3F;
                    16'h340C: data_out = 8'h40;
                    16'h340D: data_out = 8'h41;
                    16'h340E: data_out = 8'h42;
                    16'h340F: data_out = 8'h43;
                    16'h3410: data_out = 8'h44;
                    16'h3411: data_out = 8'h45;
                    16'h3412: data_out = 8'h46;
                    16'h3413: data_out = 8'h47;
                    16'h3414: data_out = 8'h48;
                    16'h3415: data_out = 8'h49;
                    16'h3416: data_out = 8'h4A;
                    16'h3417: data_out = 8'h4B;
                    16'h3418: data_out = 8'h4C;
                    16'h3419: data_out = 8'h4D;
                    16'h341A: data_out = 8'h4E;
                    16'h341B: data_out = 8'h4F;
                    16'h341C: data_out = 8'h50;
                    16'h341D: data_out = 8'h51;
                    16'h341E: data_out = 8'h52;
                    16'h341F: data_out = 8'h53;
                    16'h3420: data_out = 8'h54;
                    16'h3421: data_out = 8'h55;
                    16'h3422: data_out = 8'h56;
                    16'h3423: data_out = 8'h57;
                    16'h3424: data_out = 8'h58;
                    16'h3425: data_out = 8'h59;
                    16'h3426: data_out = 8'h5A;
                    16'h3427: data_out = 8'h5B;
                    16'h3428: data_out = 8'h5C;
                    16'h3429: data_out = 8'h5D;
                    16'h342A: data_out = 8'h5E;
                    16'h342B: data_out = 8'h5F;
                    16'h342C: data_out = 8'h60;
                    16'h342D: data_out = 8'h61;
                    16'h342E: data_out = 8'h62;
                    16'h342F: data_out = 8'h63;
                    16'h3430: data_out = 8'h64;
                    16'h3431: data_out = 8'h65;
                    16'h3432: data_out = 8'h66;
                    16'h3433: data_out = 8'h67;
                    16'h3434: data_out = 8'h68;
                    16'h3435: data_out = 8'h69;
                    16'h3436: data_out = 8'h6A;
                    16'h3437: data_out = 8'h6B;
                    16'h3438: data_out = 8'h6C;
                    16'h3439: data_out = 8'h6D;
                    16'h343A: data_out = 8'h6E;
                    16'h343B: data_out = 8'h6F;
                    16'h343C: data_out = 8'h70;
                    16'h343D: data_out = 8'h71;
                    16'h343E: data_out = 8'h72;
                    16'h343F: data_out = 8'h73;
                    16'h3440: data_out = 8'h74;
                    16'h3441: data_out = 8'h75;
                    16'h3442: data_out = 8'h76;
                    16'h3443: data_out = 8'h77;
                    16'h3444: data_out = 8'h78;
                    16'h3445: data_out = 8'h79;
                    16'h3446: data_out = 8'h7A;
                    16'h3447: data_out = 8'h7B;
                    16'h3448: data_out = 8'h7C;
                    16'h3449: data_out = 8'h7D;
                    16'h344A: data_out = 8'h7E;
                    16'h344B: data_out = 8'h7F;
                    16'h344C: data_out = 8'h80;
                    16'h344D: data_out = 8'h81;
                    16'h344E: data_out = 8'h82;
                    16'h344F: data_out = 8'h83;
                    16'h3450: data_out = 8'h84;
                    16'h3451: data_out = 8'h85;
                    16'h3452: data_out = 8'h86;
                    16'h3453: data_out = 8'h87;
                    16'h3454: data_out = 8'h88;
                    16'h3455: data_out = 8'h89;
                    16'h3456: data_out = 8'h8A;
                    16'h3457: data_out = 8'h8B;
                    16'h3458: data_out = 8'h8C;
                    16'h3459: data_out = 8'h8D;
                    16'h345A: data_out = 8'h8E;
                    16'h345B: data_out = 8'h8F;
                    16'h345C: data_out = 8'h90;
                    16'h345D: data_out = 8'h91;
                    16'h345E: data_out = 8'h92;
                    16'h345F: data_out = 8'h93;
                    16'h3460: data_out = 8'h94;
                    16'h3461: data_out = 8'h95;
                    16'h3462: data_out = 8'h96;
                    16'h3463: data_out = 8'h97;
                    16'h3464: data_out = 8'h98;
                    16'h3465: data_out = 8'h99;
                    16'h3466: data_out = 8'h9A;
                    16'h3467: data_out = 8'h9B;
                    16'h3468: data_out = 8'h9C;
                    16'h3469: data_out = 8'h9D;
                    16'h346A: data_out = 8'h9E;
                    16'h346B: data_out = 8'h9F;
                    16'h346C: data_out = 8'hA0;
                    16'h346D: data_out = 8'hA1;
                    16'h346E: data_out = 8'hA2;
                    16'h346F: data_out = 8'hA3;
                    16'h3470: data_out = 8'hA4;
                    16'h3471: data_out = 8'hA5;
                    16'h3472: data_out = 8'hA6;
                    16'h3473: data_out = 8'hA7;
                    16'h3474: data_out = 8'hA8;
                    16'h3475: data_out = 8'hA9;
                    16'h3476: data_out = 8'hAA;
                    16'h3477: data_out = 8'hAB;
                    16'h3478: data_out = 8'hAC;
                    16'h3479: data_out = 8'hAD;
                    16'h347A: data_out = 8'hAE;
                    16'h347B: data_out = 8'hAF;
                    16'h347C: data_out = 8'hB0;
                    16'h347D: data_out = 8'hB1;
                    16'h347E: data_out = 8'hB2;
                    16'h347F: data_out = 8'hB3;
                    16'h3480: data_out = 8'h34;
                    16'h3481: data_out = 8'h33;
                    16'h3482: data_out = 8'h32;
                    16'h3483: data_out = 8'h31;
                    16'h3484: data_out = 8'h30;
                    16'h3485: data_out = 8'h2F;
                    16'h3486: data_out = 8'h2E;
                    16'h3487: data_out = 8'h2D;
                    16'h3488: data_out = 8'h2C;
                    16'h3489: data_out = 8'h2B;
                    16'h348A: data_out = 8'h2A;
                    16'h348B: data_out = 8'h29;
                    16'h348C: data_out = 8'h28;
                    16'h348D: data_out = 8'h27;
                    16'h348E: data_out = 8'h26;
                    16'h348F: data_out = 8'h25;
                    16'h3490: data_out = 8'h24;
                    16'h3491: data_out = 8'h23;
                    16'h3492: data_out = 8'h22;
                    16'h3493: data_out = 8'h21;
                    16'h3494: data_out = 8'h20;
                    16'h3495: data_out = 8'h1F;
                    16'h3496: data_out = 8'h1E;
                    16'h3497: data_out = 8'h1D;
                    16'h3498: data_out = 8'h1C;
                    16'h3499: data_out = 8'h1B;
                    16'h349A: data_out = 8'h1A;
                    16'h349B: data_out = 8'h19;
                    16'h349C: data_out = 8'h18;
                    16'h349D: data_out = 8'h17;
                    16'h349E: data_out = 8'h16;
                    16'h349F: data_out = 8'h15;
                    16'h34A0: data_out = 8'h14;
                    16'h34A1: data_out = 8'h13;
                    16'h34A2: data_out = 8'h12;
                    16'h34A3: data_out = 8'h11;
                    16'h34A4: data_out = 8'h10;
                    16'h34A5: data_out = 8'hF;
                    16'h34A6: data_out = 8'hE;
                    16'h34A7: data_out = 8'hD;
                    16'h34A8: data_out = 8'hC;
                    16'h34A9: data_out = 8'hB;
                    16'h34AA: data_out = 8'hA;
                    16'h34AB: data_out = 8'h9;
                    16'h34AC: data_out = 8'h8;
                    16'h34AD: data_out = 8'h7;
                    16'h34AE: data_out = 8'h6;
                    16'h34AF: data_out = 8'h5;
                    16'h34B0: data_out = 8'h4;
                    16'h34B1: data_out = 8'h3;
                    16'h34B2: data_out = 8'h2;
                    16'h34B3: data_out = 8'h1;
                    16'h34B4: data_out = 8'h0;
                    16'h34B5: data_out = 8'h81;
                    16'h34B6: data_out = 8'h82;
                    16'h34B7: data_out = 8'h83;
                    16'h34B8: data_out = 8'h84;
                    16'h34B9: data_out = 8'h85;
                    16'h34BA: data_out = 8'h86;
                    16'h34BB: data_out = 8'h87;
                    16'h34BC: data_out = 8'h88;
                    16'h34BD: data_out = 8'h89;
                    16'h34BE: data_out = 8'h8A;
                    16'h34BF: data_out = 8'h8B;
                    16'h34C0: data_out = 8'h8C;
                    16'h34C1: data_out = 8'h8D;
                    16'h34C2: data_out = 8'h8E;
                    16'h34C3: data_out = 8'h8F;
                    16'h34C4: data_out = 8'h90;
                    16'h34C5: data_out = 8'h91;
                    16'h34C6: data_out = 8'h92;
                    16'h34C7: data_out = 8'h93;
                    16'h34C8: data_out = 8'h94;
                    16'h34C9: data_out = 8'h95;
                    16'h34CA: data_out = 8'h96;
                    16'h34CB: data_out = 8'h97;
                    16'h34CC: data_out = 8'h98;
                    16'h34CD: data_out = 8'h99;
                    16'h34CE: data_out = 8'h9A;
                    16'h34CF: data_out = 8'h9B;
                    16'h34D0: data_out = 8'h9C;
                    16'h34D1: data_out = 8'h9D;
                    16'h34D2: data_out = 8'h9E;
                    16'h34D3: data_out = 8'h9F;
                    16'h34D4: data_out = 8'hA0;
                    16'h34D5: data_out = 8'hA1;
                    16'h34D6: data_out = 8'hA2;
                    16'h34D7: data_out = 8'hA3;
                    16'h34D8: data_out = 8'hA4;
                    16'h34D9: data_out = 8'hA5;
                    16'h34DA: data_out = 8'hA6;
                    16'h34DB: data_out = 8'hA7;
                    16'h34DC: data_out = 8'hA8;
                    16'h34DD: data_out = 8'hA9;
                    16'h34DE: data_out = 8'hAA;
                    16'h34DF: data_out = 8'hAB;
                    16'h34E0: data_out = 8'hAC;
                    16'h34E1: data_out = 8'hAD;
                    16'h34E2: data_out = 8'hAE;
                    16'h34E3: data_out = 8'hAF;
                    16'h34E4: data_out = 8'hB0;
                    16'h34E5: data_out = 8'hB1;
                    16'h34E6: data_out = 8'hB2;
                    16'h34E7: data_out = 8'hB3;
                    16'h34E8: data_out = 8'hB4;
                    16'h34E9: data_out = 8'hB5;
                    16'h34EA: data_out = 8'hB6;
                    16'h34EB: data_out = 8'hB7;
                    16'h34EC: data_out = 8'hB8;
                    16'h34ED: data_out = 8'hB9;
                    16'h34EE: data_out = 8'hBA;
                    16'h34EF: data_out = 8'hBB;
                    16'h34F0: data_out = 8'hBC;
                    16'h34F1: data_out = 8'hBD;
                    16'h34F2: data_out = 8'hBE;
                    16'h34F3: data_out = 8'hBF;
                    16'h34F4: data_out = 8'hC0;
                    16'h34F5: data_out = 8'hC1;
                    16'h34F6: data_out = 8'hC2;
                    16'h34F7: data_out = 8'hC3;
                    16'h34F8: data_out = 8'hC4;
                    16'h34F9: data_out = 8'hC5;
                    16'h34FA: data_out = 8'hC6;
                    16'h34FB: data_out = 8'hC7;
                    16'h34FC: data_out = 8'hC8;
                    16'h34FD: data_out = 8'hC9;
                    16'h34FE: data_out = 8'hCA;
                    16'h34FF: data_out = 8'hCB;
                    16'h3500: data_out = 8'h35;
                    16'h3501: data_out = 8'h36;
                    16'h3502: data_out = 8'h37;
                    16'h3503: data_out = 8'h38;
                    16'h3504: data_out = 8'h39;
                    16'h3505: data_out = 8'h3A;
                    16'h3506: data_out = 8'h3B;
                    16'h3507: data_out = 8'h3C;
                    16'h3508: data_out = 8'h3D;
                    16'h3509: data_out = 8'h3E;
                    16'h350A: data_out = 8'h3F;
                    16'h350B: data_out = 8'h40;
                    16'h350C: data_out = 8'h41;
                    16'h350D: data_out = 8'h42;
                    16'h350E: data_out = 8'h43;
                    16'h350F: data_out = 8'h44;
                    16'h3510: data_out = 8'h45;
                    16'h3511: data_out = 8'h46;
                    16'h3512: data_out = 8'h47;
                    16'h3513: data_out = 8'h48;
                    16'h3514: data_out = 8'h49;
                    16'h3515: data_out = 8'h4A;
                    16'h3516: data_out = 8'h4B;
                    16'h3517: data_out = 8'h4C;
                    16'h3518: data_out = 8'h4D;
                    16'h3519: data_out = 8'h4E;
                    16'h351A: data_out = 8'h4F;
                    16'h351B: data_out = 8'h50;
                    16'h351C: data_out = 8'h51;
                    16'h351D: data_out = 8'h52;
                    16'h351E: data_out = 8'h53;
                    16'h351F: data_out = 8'h54;
                    16'h3520: data_out = 8'h55;
                    16'h3521: data_out = 8'h56;
                    16'h3522: data_out = 8'h57;
                    16'h3523: data_out = 8'h58;
                    16'h3524: data_out = 8'h59;
                    16'h3525: data_out = 8'h5A;
                    16'h3526: data_out = 8'h5B;
                    16'h3527: data_out = 8'h5C;
                    16'h3528: data_out = 8'h5D;
                    16'h3529: data_out = 8'h5E;
                    16'h352A: data_out = 8'h5F;
                    16'h352B: data_out = 8'h60;
                    16'h352C: data_out = 8'h61;
                    16'h352D: data_out = 8'h62;
                    16'h352E: data_out = 8'h63;
                    16'h352F: data_out = 8'h64;
                    16'h3530: data_out = 8'h65;
                    16'h3531: data_out = 8'h66;
                    16'h3532: data_out = 8'h67;
                    16'h3533: data_out = 8'h68;
                    16'h3534: data_out = 8'h69;
                    16'h3535: data_out = 8'h6A;
                    16'h3536: data_out = 8'h6B;
                    16'h3537: data_out = 8'h6C;
                    16'h3538: data_out = 8'h6D;
                    16'h3539: data_out = 8'h6E;
                    16'h353A: data_out = 8'h6F;
                    16'h353B: data_out = 8'h70;
                    16'h353C: data_out = 8'h71;
                    16'h353D: data_out = 8'h72;
                    16'h353E: data_out = 8'h73;
                    16'h353F: data_out = 8'h74;
                    16'h3540: data_out = 8'h75;
                    16'h3541: data_out = 8'h76;
                    16'h3542: data_out = 8'h77;
                    16'h3543: data_out = 8'h78;
                    16'h3544: data_out = 8'h79;
                    16'h3545: data_out = 8'h7A;
                    16'h3546: data_out = 8'h7B;
                    16'h3547: data_out = 8'h7C;
                    16'h3548: data_out = 8'h7D;
                    16'h3549: data_out = 8'h7E;
                    16'h354A: data_out = 8'h7F;
                    16'h354B: data_out = 8'h80;
                    16'h354C: data_out = 8'h81;
                    16'h354D: data_out = 8'h82;
                    16'h354E: data_out = 8'h83;
                    16'h354F: data_out = 8'h84;
                    16'h3550: data_out = 8'h85;
                    16'h3551: data_out = 8'h86;
                    16'h3552: data_out = 8'h87;
                    16'h3553: data_out = 8'h88;
                    16'h3554: data_out = 8'h89;
                    16'h3555: data_out = 8'h8A;
                    16'h3556: data_out = 8'h8B;
                    16'h3557: data_out = 8'h8C;
                    16'h3558: data_out = 8'h8D;
                    16'h3559: data_out = 8'h8E;
                    16'h355A: data_out = 8'h8F;
                    16'h355B: data_out = 8'h90;
                    16'h355C: data_out = 8'h91;
                    16'h355D: data_out = 8'h92;
                    16'h355E: data_out = 8'h93;
                    16'h355F: data_out = 8'h94;
                    16'h3560: data_out = 8'h95;
                    16'h3561: data_out = 8'h96;
                    16'h3562: data_out = 8'h97;
                    16'h3563: data_out = 8'h98;
                    16'h3564: data_out = 8'h99;
                    16'h3565: data_out = 8'h9A;
                    16'h3566: data_out = 8'h9B;
                    16'h3567: data_out = 8'h9C;
                    16'h3568: data_out = 8'h9D;
                    16'h3569: data_out = 8'h9E;
                    16'h356A: data_out = 8'h9F;
                    16'h356B: data_out = 8'hA0;
                    16'h356C: data_out = 8'hA1;
                    16'h356D: data_out = 8'hA2;
                    16'h356E: data_out = 8'hA3;
                    16'h356F: data_out = 8'hA4;
                    16'h3570: data_out = 8'hA5;
                    16'h3571: data_out = 8'hA6;
                    16'h3572: data_out = 8'hA7;
                    16'h3573: data_out = 8'hA8;
                    16'h3574: data_out = 8'hA9;
                    16'h3575: data_out = 8'hAA;
                    16'h3576: data_out = 8'hAB;
                    16'h3577: data_out = 8'hAC;
                    16'h3578: data_out = 8'hAD;
                    16'h3579: data_out = 8'hAE;
                    16'h357A: data_out = 8'hAF;
                    16'h357B: data_out = 8'hB0;
                    16'h357C: data_out = 8'hB1;
                    16'h357D: data_out = 8'hB2;
                    16'h357E: data_out = 8'hB3;
                    16'h357F: data_out = 8'hB4;
                    16'h3580: data_out = 8'h35;
                    16'h3581: data_out = 8'h34;
                    16'h3582: data_out = 8'h33;
                    16'h3583: data_out = 8'h32;
                    16'h3584: data_out = 8'h31;
                    16'h3585: data_out = 8'h30;
                    16'h3586: data_out = 8'h2F;
                    16'h3587: data_out = 8'h2E;
                    16'h3588: data_out = 8'h2D;
                    16'h3589: data_out = 8'h2C;
                    16'h358A: data_out = 8'h2B;
                    16'h358B: data_out = 8'h2A;
                    16'h358C: data_out = 8'h29;
                    16'h358D: data_out = 8'h28;
                    16'h358E: data_out = 8'h27;
                    16'h358F: data_out = 8'h26;
                    16'h3590: data_out = 8'h25;
                    16'h3591: data_out = 8'h24;
                    16'h3592: data_out = 8'h23;
                    16'h3593: data_out = 8'h22;
                    16'h3594: data_out = 8'h21;
                    16'h3595: data_out = 8'h20;
                    16'h3596: data_out = 8'h1F;
                    16'h3597: data_out = 8'h1E;
                    16'h3598: data_out = 8'h1D;
                    16'h3599: data_out = 8'h1C;
                    16'h359A: data_out = 8'h1B;
                    16'h359B: data_out = 8'h1A;
                    16'h359C: data_out = 8'h19;
                    16'h359D: data_out = 8'h18;
                    16'h359E: data_out = 8'h17;
                    16'h359F: data_out = 8'h16;
                    16'h35A0: data_out = 8'h15;
                    16'h35A1: data_out = 8'h14;
                    16'h35A2: data_out = 8'h13;
                    16'h35A3: data_out = 8'h12;
                    16'h35A4: data_out = 8'h11;
                    16'h35A5: data_out = 8'h10;
                    16'h35A6: data_out = 8'hF;
                    16'h35A7: data_out = 8'hE;
                    16'h35A8: data_out = 8'hD;
                    16'h35A9: data_out = 8'hC;
                    16'h35AA: data_out = 8'hB;
                    16'h35AB: data_out = 8'hA;
                    16'h35AC: data_out = 8'h9;
                    16'h35AD: data_out = 8'h8;
                    16'h35AE: data_out = 8'h7;
                    16'h35AF: data_out = 8'h6;
                    16'h35B0: data_out = 8'h5;
                    16'h35B1: data_out = 8'h4;
                    16'h35B2: data_out = 8'h3;
                    16'h35B3: data_out = 8'h2;
                    16'h35B4: data_out = 8'h1;
                    16'h35B5: data_out = 8'h0;
                    16'h35B6: data_out = 8'h81;
                    16'h35B7: data_out = 8'h82;
                    16'h35B8: data_out = 8'h83;
                    16'h35B9: data_out = 8'h84;
                    16'h35BA: data_out = 8'h85;
                    16'h35BB: data_out = 8'h86;
                    16'h35BC: data_out = 8'h87;
                    16'h35BD: data_out = 8'h88;
                    16'h35BE: data_out = 8'h89;
                    16'h35BF: data_out = 8'h8A;
                    16'h35C0: data_out = 8'h8B;
                    16'h35C1: data_out = 8'h8C;
                    16'h35C2: data_out = 8'h8D;
                    16'h35C3: data_out = 8'h8E;
                    16'h35C4: data_out = 8'h8F;
                    16'h35C5: data_out = 8'h90;
                    16'h35C6: data_out = 8'h91;
                    16'h35C7: data_out = 8'h92;
                    16'h35C8: data_out = 8'h93;
                    16'h35C9: data_out = 8'h94;
                    16'h35CA: data_out = 8'h95;
                    16'h35CB: data_out = 8'h96;
                    16'h35CC: data_out = 8'h97;
                    16'h35CD: data_out = 8'h98;
                    16'h35CE: data_out = 8'h99;
                    16'h35CF: data_out = 8'h9A;
                    16'h35D0: data_out = 8'h9B;
                    16'h35D1: data_out = 8'h9C;
                    16'h35D2: data_out = 8'h9D;
                    16'h35D3: data_out = 8'h9E;
                    16'h35D4: data_out = 8'h9F;
                    16'h35D5: data_out = 8'hA0;
                    16'h35D6: data_out = 8'hA1;
                    16'h35D7: data_out = 8'hA2;
                    16'h35D8: data_out = 8'hA3;
                    16'h35D9: data_out = 8'hA4;
                    16'h35DA: data_out = 8'hA5;
                    16'h35DB: data_out = 8'hA6;
                    16'h35DC: data_out = 8'hA7;
                    16'h35DD: data_out = 8'hA8;
                    16'h35DE: data_out = 8'hA9;
                    16'h35DF: data_out = 8'hAA;
                    16'h35E0: data_out = 8'hAB;
                    16'h35E1: data_out = 8'hAC;
                    16'h35E2: data_out = 8'hAD;
                    16'h35E3: data_out = 8'hAE;
                    16'h35E4: data_out = 8'hAF;
                    16'h35E5: data_out = 8'hB0;
                    16'h35E6: data_out = 8'hB1;
                    16'h35E7: data_out = 8'hB2;
                    16'h35E8: data_out = 8'hB3;
                    16'h35E9: data_out = 8'hB4;
                    16'h35EA: data_out = 8'hB5;
                    16'h35EB: data_out = 8'hB6;
                    16'h35EC: data_out = 8'hB7;
                    16'h35ED: data_out = 8'hB8;
                    16'h35EE: data_out = 8'hB9;
                    16'h35EF: data_out = 8'hBA;
                    16'h35F0: data_out = 8'hBB;
                    16'h35F1: data_out = 8'hBC;
                    16'h35F2: data_out = 8'hBD;
                    16'h35F3: data_out = 8'hBE;
                    16'h35F4: data_out = 8'hBF;
                    16'h35F5: data_out = 8'hC0;
                    16'h35F6: data_out = 8'hC1;
                    16'h35F7: data_out = 8'hC2;
                    16'h35F8: data_out = 8'hC3;
                    16'h35F9: data_out = 8'hC4;
                    16'h35FA: data_out = 8'hC5;
                    16'h35FB: data_out = 8'hC6;
                    16'h35FC: data_out = 8'hC7;
                    16'h35FD: data_out = 8'hC8;
                    16'h35FE: data_out = 8'hC9;
                    16'h35FF: data_out = 8'hCA;
                    16'h3600: data_out = 8'h36;
                    16'h3601: data_out = 8'h37;
                    16'h3602: data_out = 8'h38;
                    16'h3603: data_out = 8'h39;
                    16'h3604: data_out = 8'h3A;
                    16'h3605: data_out = 8'h3B;
                    16'h3606: data_out = 8'h3C;
                    16'h3607: data_out = 8'h3D;
                    16'h3608: data_out = 8'h3E;
                    16'h3609: data_out = 8'h3F;
                    16'h360A: data_out = 8'h40;
                    16'h360B: data_out = 8'h41;
                    16'h360C: data_out = 8'h42;
                    16'h360D: data_out = 8'h43;
                    16'h360E: data_out = 8'h44;
                    16'h360F: data_out = 8'h45;
                    16'h3610: data_out = 8'h46;
                    16'h3611: data_out = 8'h47;
                    16'h3612: data_out = 8'h48;
                    16'h3613: data_out = 8'h49;
                    16'h3614: data_out = 8'h4A;
                    16'h3615: data_out = 8'h4B;
                    16'h3616: data_out = 8'h4C;
                    16'h3617: data_out = 8'h4D;
                    16'h3618: data_out = 8'h4E;
                    16'h3619: data_out = 8'h4F;
                    16'h361A: data_out = 8'h50;
                    16'h361B: data_out = 8'h51;
                    16'h361C: data_out = 8'h52;
                    16'h361D: data_out = 8'h53;
                    16'h361E: data_out = 8'h54;
                    16'h361F: data_out = 8'h55;
                    16'h3620: data_out = 8'h56;
                    16'h3621: data_out = 8'h57;
                    16'h3622: data_out = 8'h58;
                    16'h3623: data_out = 8'h59;
                    16'h3624: data_out = 8'h5A;
                    16'h3625: data_out = 8'h5B;
                    16'h3626: data_out = 8'h5C;
                    16'h3627: data_out = 8'h5D;
                    16'h3628: data_out = 8'h5E;
                    16'h3629: data_out = 8'h5F;
                    16'h362A: data_out = 8'h60;
                    16'h362B: data_out = 8'h61;
                    16'h362C: data_out = 8'h62;
                    16'h362D: data_out = 8'h63;
                    16'h362E: data_out = 8'h64;
                    16'h362F: data_out = 8'h65;
                    16'h3630: data_out = 8'h66;
                    16'h3631: data_out = 8'h67;
                    16'h3632: data_out = 8'h68;
                    16'h3633: data_out = 8'h69;
                    16'h3634: data_out = 8'h6A;
                    16'h3635: data_out = 8'h6B;
                    16'h3636: data_out = 8'h6C;
                    16'h3637: data_out = 8'h6D;
                    16'h3638: data_out = 8'h6E;
                    16'h3639: data_out = 8'h6F;
                    16'h363A: data_out = 8'h70;
                    16'h363B: data_out = 8'h71;
                    16'h363C: data_out = 8'h72;
                    16'h363D: data_out = 8'h73;
                    16'h363E: data_out = 8'h74;
                    16'h363F: data_out = 8'h75;
                    16'h3640: data_out = 8'h76;
                    16'h3641: data_out = 8'h77;
                    16'h3642: data_out = 8'h78;
                    16'h3643: data_out = 8'h79;
                    16'h3644: data_out = 8'h7A;
                    16'h3645: data_out = 8'h7B;
                    16'h3646: data_out = 8'h7C;
                    16'h3647: data_out = 8'h7D;
                    16'h3648: data_out = 8'h7E;
                    16'h3649: data_out = 8'h7F;
                    16'h364A: data_out = 8'h80;
                    16'h364B: data_out = 8'h81;
                    16'h364C: data_out = 8'h82;
                    16'h364D: data_out = 8'h83;
                    16'h364E: data_out = 8'h84;
                    16'h364F: data_out = 8'h85;
                    16'h3650: data_out = 8'h86;
                    16'h3651: data_out = 8'h87;
                    16'h3652: data_out = 8'h88;
                    16'h3653: data_out = 8'h89;
                    16'h3654: data_out = 8'h8A;
                    16'h3655: data_out = 8'h8B;
                    16'h3656: data_out = 8'h8C;
                    16'h3657: data_out = 8'h8D;
                    16'h3658: data_out = 8'h8E;
                    16'h3659: data_out = 8'h8F;
                    16'h365A: data_out = 8'h90;
                    16'h365B: data_out = 8'h91;
                    16'h365C: data_out = 8'h92;
                    16'h365D: data_out = 8'h93;
                    16'h365E: data_out = 8'h94;
                    16'h365F: data_out = 8'h95;
                    16'h3660: data_out = 8'h96;
                    16'h3661: data_out = 8'h97;
                    16'h3662: data_out = 8'h98;
                    16'h3663: data_out = 8'h99;
                    16'h3664: data_out = 8'h9A;
                    16'h3665: data_out = 8'h9B;
                    16'h3666: data_out = 8'h9C;
                    16'h3667: data_out = 8'h9D;
                    16'h3668: data_out = 8'h9E;
                    16'h3669: data_out = 8'h9F;
                    16'h366A: data_out = 8'hA0;
                    16'h366B: data_out = 8'hA1;
                    16'h366C: data_out = 8'hA2;
                    16'h366D: data_out = 8'hA3;
                    16'h366E: data_out = 8'hA4;
                    16'h366F: data_out = 8'hA5;
                    16'h3670: data_out = 8'hA6;
                    16'h3671: data_out = 8'hA7;
                    16'h3672: data_out = 8'hA8;
                    16'h3673: data_out = 8'hA9;
                    16'h3674: data_out = 8'hAA;
                    16'h3675: data_out = 8'hAB;
                    16'h3676: data_out = 8'hAC;
                    16'h3677: data_out = 8'hAD;
                    16'h3678: data_out = 8'hAE;
                    16'h3679: data_out = 8'hAF;
                    16'h367A: data_out = 8'hB0;
                    16'h367B: data_out = 8'hB1;
                    16'h367C: data_out = 8'hB2;
                    16'h367D: data_out = 8'hB3;
                    16'h367E: data_out = 8'hB4;
                    16'h367F: data_out = 8'hB5;
                    16'h3680: data_out = 8'h36;
                    16'h3681: data_out = 8'h35;
                    16'h3682: data_out = 8'h34;
                    16'h3683: data_out = 8'h33;
                    16'h3684: data_out = 8'h32;
                    16'h3685: data_out = 8'h31;
                    16'h3686: data_out = 8'h30;
                    16'h3687: data_out = 8'h2F;
                    16'h3688: data_out = 8'h2E;
                    16'h3689: data_out = 8'h2D;
                    16'h368A: data_out = 8'h2C;
                    16'h368B: data_out = 8'h2B;
                    16'h368C: data_out = 8'h2A;
                    16'h368D: data_out = 8'h29;
                    16'h368E: data_out = 8'h28;
                    16'h368F: data_out = 8'h27;
                    16'h3690: data_out = 8'h26;
                    16'h3691: data_out = 8'h25;
                    16'h3692: data_out = 8'h24;
                    16'h3693: data_out = 8'h23;
                    16'h3694: data_out = 8'h22;
                    16'h3695: data_out = 8'h21;
                    16'h3696: data_out = 8'h20;
                    16'h3697: data_out = 8'h1F;
                    16'h3698: data_out = 8'h1E;
                    16'h3699: data_out = 8'h1D;
                    16'h369A: data_out = 8'h1C;
                    16'h369B: data_out = 8'h1B;
                    16'h369C: data_out = 8'h1A;
                    16'h369D: data_out = 8'h19;
                    16'h369E: data_out = 8'h18;
                    16'h369F: data_out = 8'h17;
                    16'h36A0: data_out = 8'h16;
                    16'h36A1: data_out = 8'h15;
                    16'h36A2: data_out = 8'h14;
                    16'h36A3: data_out = 8'h13;
                    16'h36A4: data_out = 8'h12;
                    16'h36A5: data_out = 8'h11;
                    16'h36A6: data_out = 8'h10;
                    16'h36A7: data_out = 8'hF;
                    16'h36A8: data_out = 8'hE;
                    16'h36A9: data_out = 8'hD;
                    16'h36AA: data_out = 8'hC;
                    16'h36AB: data_out = 8'hB;
                    16'h36AC: data_out = 8'hA;
                    16'h36AD: data_out = 8'h9;
                    16'h36AE: data_out = 8'h8;
                    16'h36AF: data_out = 8'h7;
                    16'h36B0: data_out = 8'h6;
                    16'h36B1: data_out = 8'h5;
                    16'h36B2: data_out = 8'h4;
                    16'h36B3: data_out = 8'h3;
                    16'h36B4: data_out = 8'h2;
                    16'h36B5: data_out = 8'h1;
                    16'h36B6: data_out = 8'h0;
                    16'h36B7: data_out = 8'h81;
                    16'h36B8: data_out = 8'h82;
                    16'h36B9: data_out = 8'h83;
                    16'h36BA: data_out = 8'h84;
                    16'h36BB: data_out = 8'h85;
                    16'h36BC: data_out = 8'h86;
                    16'h36BD: data_out = 8'h87;
                    16'h36BE: data_out = 8'h88;
                    16'h36BF: data_out = 8'h89;
                    16'h36C0: data_out = 8'h8A;
                    16'h36C1: data_out = 8'h8B;
                    16'h36C2: data_out = 8'h8C;
                    16'h36C3: data_out = 8'h8D;
                    16'h36C4: data_out = 8'h8E;
                    16'h36C5: data_out = 8'h8F;
                    16'h36C6: data_out = 8'h90;
                    16'h36C7: data_out = 8'h91;
                    16'h36C8: data_out = 8'h92;
                    16'h36C9: data_out = 8'h93;
                    16'h36CA: data_out = 8'h94;
                    16'h36CB: data_out = 8'h95;
                    16'h36CC: data_out = 8'h96;
                    16'h36CD: data_out = 8'h97;
                    16'h36CE: data_out = 8'h98;
                    16'h36CF: data_out = 8'h99;
                    16'h36D0: data_out = 8'h9A;
                    16'h36D1: data_out = 8'h9B;
                    16'h36D2: data_out = 8'h9C;
                    16'h36D3: data_out = 8'h9D;
                    16'h36D4: data_out = 8'h9E;
                    16'h36D5: data_out = 8'h9F;
                    16'h36D6: data_out = 8'hA0;
                    16'h36D7: data_out = 8'hA1;
                    16'h36D8: data_out = 8'hA2;
                    16'h36D9: data_out = 8'hA3;
                    16'h36DA: data_out = 8'hA4;
                    16'h36DB: data_out = 8'hA5;
                    16'h36DC: data_out = 8'hA6;
                    16'h36DD: data_out = 8'hA7;
                    16'h36DE: data_out = 8'hA8;
                    16'h36DF: data_out = 8'hA9;
                    16'h36E0: data_out = 8'hAA;
                    16'h36E1: data_out = 8'hAB;
                    16'h36E2: data_out = 8'hAC;
                    16'h36E3: data_out = 8'hAD;
                    16'h36E4: data_out = 8'hAE;
                    16'h36E5: data_out = 8'hAF;
                    16'h36E6: data_out = 8'hB0;
                    16'h36E7: data_out = 8'hB1;
                    16'h36E8: data_out = 8'hB2;
                    16'h36E9: data_out = 8'hB3;
                    16'h36EA: data_out = 8'hB4;
                    16'h36EB: data_out = 8'hB5;
                    16'h36EC: data_out = 8'hB6;
                    16'h36ED: data_out = 8'hB7;
                    16'h36EE: data_out = 8'hB8;
                    16'h36EF: data_out = 8'hB9;
                    16'h36F0: data_out = 8'hBA;
                    16'h36F1: data_out = 8'hBB;
                    16'h36F2: data_out = 8'hBC;
                    16'h36F3: data_out = 8'hBD;
                    16'h36F4: data_out = 8'hBE;
                    16'h36F5: data_out = 8'hBF;
                    16'h36F6: data_out = 8'hC0;
                    16'h36F7: data_out = 8'hC1;
                    16'h36F8: data_out = 8'hC2;
                    16'h36F9: data_out = 8'hC3;
                    16'h36FA: data_out = 8'hC4;
                    16'h36FB: data_out = 8'hC5;
                    16'h36FC: data_out = 8'hC6;
                    16'h36FD: data_out = 8'hC7;
                    16'h36FE: data_out = 8'hC8;
                    16'h36FF: data_out = 8'hC9;
                    16'h3700: data_out = 8'h37;
                    16'h3701: data_out = 8'h38;
                    16'h3702: data_out = 8'h39;
                    16'h3703: data_out = 8'h3A;
                    16'h3704: data_out = 8'h3B;
                    16'h3705: data_out = 8'h3C;
                    16'h3706: data_out = 8'h3D;
                    16'h3707: data_out = 8'h3E;
                    16'h3708: data_out = 8'h3F;
                    16'h3709: data_out = 8'h40;
                    16'h370A: data_out = 8'h41;
                    16'h370B: data_out = 8'h42;
                    16'h370C: data_out = 8'h43;
                    16'h370D: data_out = 8'h44;
                    16'h370E: data_out = 8'h45;
                    16'h370F: data_out = 8'h46;
                    16'h3710: data_out = 8'h47;
                    16'h3711: data_out = 8'h48;
                    16'h3712: data_out = 8'h49;
                    16'h3713: data_out = 8'h4A;
                    16'h3714: data_out = 8'h4B;
                    16'h3715: data_out = 8'h4C;
                    16'h3716: data_out = 8'h4D;
                    16'h3717: data_out = 8'h4E;
                    16'h3718: data_out = 8'h4F;
                    16'h3719: data_out = 8'h50;
                    16'h371A: data_out = 8'h51;
                    16'h371B: data_out = 8'h52;
                    16'h371C: data_out = 8'h53;
                    16'h371D: data_out = 8'h54;
                    16'h371E: data_out = 8'h55;
                    16'h371F: data_out = 8'h56;
                    16'h3720: data_out = 8'h57;
                    16'h3721: data_out = 8'h58;
                    16'h3722: data_out = 8'h59;
                    16'h3723: data_out = 8'h5A;
                    16'h3724: data_out = 8'h5B;
                    16'h3725: data_out = 8'h5C;
                    16'h3726: data_out = 8'h5D;
                    16'h3727: data_out = 8'h5E;
                    16'h3728: data_out = 8'h5F;
                    16'h3729: data_out = 8'h60;
                    16'h372A: data_out = 8'h61;
                    16'h372B: data_out = 8'h62;
                    16'h372C: data_out = 8'h63;
                    16'h372D: data_out = 8'h64;
                    16'h372E: data_out = 8'h65;
                    16'h372F: data_out = 8'h66;
                    16'h3730: data_out = 8'h67;
                    16'h3731: data_out = 8'h68;
                    16'h3732: data_out = 8'h69;
                    16'h3733: data_out = 8'h6A;
                    16'h3734: data_out = 8'h6B;
                    16'h3735: data_out = 8'h6C;
                    16'h3736: data_out = 8'h6D;
                    16'h3737: data_out = 8'h6E;
                    16'h3738: data_out = 8'h6F;
                    16'h3739: data_out = 8'h70;
                    16'h373A: data_out = 8'h71;
                    16'h373B: data_out = 8'h72;
                    16'h373C: data_out = 8'h73;
                    16'h373D: data_out = 8'h74;
                    16'h373E: data_out = 8'h75;
                    16'h373F: data_out = 8'h76;
                    16'h3740: data_out = 8'h77;
                    16'h3741: data_out = 8'h78;
                    16'h3742: data_out = 8'h79;
                    16'h3743: data_out = 8'h7A;
                    16'h3744: data_out = 8'h7B;
                    16'h3745: data_out = 8'h7C;
                    16'h3746: data_out = 8'h7D;
                    16'h3747: data_out = 8'h7E;
                    16'h3748: data_out = 8'h7F;
                    16'h3749: data_out = 8'h80;
                    16'h374A: data_out = 8'h81;
                    16'h374B: data_out = 8'h82;
                    16'h374C: data_out = 8'h83;
                    16'h374D: data_out = 8'h84;
                    16'h374E: data_out = 8'h85;
                    16'h374F: data_out = 8'h86;
                    16'h3750: data_out = 8'h87;
                    16'h3751: data_out = 8'h88;
                    16'h3752: data_out = 8'h89;
                    16'h3753: data_out = 8'h8A;
                    16'h3754: data_out = 8'h8B;
                    16'h3755: data_out = 8'h8C;
                    16'h3756: data_out = 8'h8D;
                    16'h3757: data_out = 8'h8E;
                    16'h3758: data_out = 8'h8F;
                    16'h3759: data_out = 8'h90;
                    16'h375A: data_out = 8'h91;
                    16'h375B: data_out = 8'h92;
                    16'h375C: data_out = 8'h93;
                    16'h375D: data_out = 8'h94;
                    16'h375E: data_out = 8'h95;
                    16'h375F: data_out = 8'h96;
                    16'h3760: data_out = 8'h97;
                    16'h3761: data_out = 8'h98;
                    16'h3762: data_out = 8'h99;
                    16'h3763: data_out = 8'h9A;
                    16'h3764: data_out = 8'h9B;
                    16'h3765: data_out = 8'h9C;
                    16'h3766: data_out = 8'h9D;
                    16'h3767: data_out = 8'h9E;
                    16'h3768: data_out = 8'h9F;
                    16'h3769: data_out = 8'hA0;
                    16'h376A: data_out = 8'hA1;
                    16'h376B: data_out = 8'hA2;
                    16'h376C: data_out = 8'hA3;
                    16'h376D: data_out = 8'hA4;
                    16'h376E: data_out = 8'hA5;
                    16'h376F: data_out = 8'hA6;
                    16'h3770: data_out = 8'hA7;
                    16'h3771: data_out = 8'hA8;
                    16'h3772: data_out = 8'hA9;
                    16'h3773: data_out = 8'hAA;
                    16'h3774: data_out = 8'hAB;
                    16'h3775: data_out = 8'hAC;
                    16'h3776: data_out = 8'hAD;
                    16'h3777: data_out = 8'hAE;
                    16'h3778: data_out = 8'hAF;
                    16'h3779: data_out = 8'hB0;
                    16'h377A: data_out = 8'hB1;
                    16'h377B: data_out = 8'hB2;
                    16'h377C: data_out = 8'hB3;
                    16'h377D: data_out = 8'hB4;
                    16'h377E: data_out = 8'hB5;
                    16'h377F: data_out = 8'hB6;
                    16'h3780: data_out = 8'h37;
                    16'h3781: data_out = 8'h36;
                    16'h3782: data_out = 8'h35;
                    16'h3783: data_out = 8'h34;
                    16'h3784: data_out = 8'h33;
                    16'h3785: data_out = 8'h32;
                    16'h3786: data_out = 8'h31;
                    16'h3787: data_out = 8'h30;
                    16'h3788: data_out = 8'h2F;
                    16'h3789: data_out = 8'h2E;
                    16'h378A: data_out = 8'h2D;
                    16'h378B: data_out = 8'h2C;
                    16'h378C: data_out = 8'h2B;
                    16'h378D: data_out = 8'h2A;
                    16'h378E: data_out = 8'h29;
                    16'h378F: data_out = 8'h28;
                    16'h3790: data_out = 8'h27;
                    16'h3791: data_out = 8'h26;
                    16'h3792: data_out = 8'h25;
                    16'h3793: data_out = 8'h24;
                    16'h3794: data_out = 8'h23;
                    16'h3795: data_out = 8'h22;
                    16'h3796: data_out = 8'h21;
                    16'h3797: data_out = 8'h20;
                    16'h3798: data_out = 8'h1F;
                    16'h3799: data_out = 8'h1E;
                    16'h379A: data_out = 8'h1D;
                    16'h379B: data_out = 8'h1C;
                    16'h379C: data_out = 8'h1B;
                    16'h379D: data_out = 8'h1A;
                    16'h379E: data_out = 8'h19;
                    16'h379F: data_out = 8'h18;
                    16'h37A0: data_out = 8'h17;
                    16'h37A1: data_out = 8'h16;
                    16'h37A2: data_out = 8'h15;
                    16'h37A3: data_out = 8'h14;
                    16'h37A4: data_out = 8'h13;
                    16'h37A5: data_out = 8'h12;
                    16'h37A6: data_out = 8'h11;
                    16'h37A7: data_out = 8'h10;
                    16'h37A8: data_out = 8'hF;
                    16'h37A9: data_out = 8'hE;
                    16'h37AA: data_out = 8'hD;
                    16'h37AB: data_out = 8'hC;
                    16'h37AC: data_out = 8'hB;
                    16'h37AD: data_out = 8'hA;
                    16'h37AE: data_out = 8'h9;
                    16'h37AF: data_out = 8'h8;
                    16'h37B0: data_out = 8'h7;
                    16'h37B1: data_out = 8'h6;
                    16'h37B2: data_out = 8'h5;
                    16'h37B3: data_out = 8'h4;
                    16'h37B4: data_out = 8'h3;
                    16'h37B5: data_out = 8'h2;
                    16'h37B6: data_out = 8'h1;
                    16'h37B7: data_out = 8'h0;
                    16'h37B8: data_out = 8'h81;
                    16'h37B9: data_out = 8'h82;
                    16'h37BA: data_out = 8'h83;
                    16'h37BB: data_out = 8'h84;
                    16'h37BC: data_out = 8'h85;
                    16'h37BD: data_out = 8'h86;
                    16'h37BE: data_out = 8'h87;
                    16'h37BF: data_out = 8'h88;
                    16'h37C0: data_out = 8'h89;
                    16'h37C1: data_out = 8'h8A;
                    16'h37C2: data_out = 8'h8B;
                    16'h37C3: data_out = 8'h8C;
                    16'h37C4: data_out = 8'h8D;
                    16'h37C5: data_out = 8'h8E;
                    16'h37C6: data_out = 8'h8F;
                    16'h37C7: data_out = 8'h90;
                    16'h37C8: data_out = 8'h91;
                    16'h37C9: data_out = 8'h92;
                    16'h37CA: data_out = 8'h93;
                    16'h37CB: data_out = 8'h94;
                    16'h37CC: data_out = 8'h95;
                    16'h37CD: data_out = 8'h96;
                    16'h37CE: data_out = 8'h97;
                    16'h37CF: data_out = 8'h98;
                    16'h37D0: data_out = 8'h99;
                    16'h37D1: data_out = 8'h9A;
                    16'h37D2: data_out = 8'h9B;
                    16'h37D3: data_out = 8'h9C;
                    16'h37D4: data_out = 8'h9D;
                    16'h37D5: data_out = 8'h9E;
                    16'h37D6: data_out = 8'h9F;
                    16'h37D7: data_out = 8'hA0;
                    16'h37D8: data_out = 8'hA1;
                    16'h37D9: data_out = 8'hA2;
                    16'h37DA: data_out = 8'hA3;
                    16'h37DB: data_out = 8'hA4;
                    16'h37DC: data_out = 8'hA5;
                    16'h37DD: data_out = 8'hA6;
                    16'h37DE: data_out = 8'hA7;
                    16'h37DF: data_out = 8'hA8;
                    16'h37E0: data_out = 8'hA9;
                    16'h37E1: data_out = 8'hAA;
                    16'h37E2: data_out = 8'hAB;
                    16'h37E3: data_out = 8'hAC;
                    16'h37E4: data_out = 8'hAD;
                    16'h37E5: data_out = 8'hAE;
                    16'h37E6: data_out = 8'hAF;
                    16'h37E7: data_out = 8'hB0;
                    16'h37E8: data_out = 8'hB1;
                    16'h37E9: data_out = 8'hB2;
                    16'h37EA: data_out = 8'hB3;
                    16'h37EB: data_out = 8'hB4;
                    16'h37EC: data_out = 8'hB5;
                    16'h37ED: data_out = 8'hB6;
                    16'h37EE: data_out = 8'hB7;
                    16'h37EF: data_out = 8'hB8;
                    16'h37F0: data_out = 8'hB9;
                    16'h37F1: data_out = 8'hBA;
                    16'h37F2: data_out = 8'hBB;
                    16'h37F3: data_out = 8'hBC;
                    16'h37F4: data_out = 8'hBD;
                    16'h37F5: data_out = 8'hBE;
                    16'h37F6: data_out = 8'hBF;
                    16'h37F7: data_out = 8'hC0;
                    16'h37F8: data_out = 8'hC1;
                    16'h37F9: data_out = 8'hC2;
                    16'h37FA: data_out = 8'hC3;
                    16'h37FB: data_out = 8'hC4;
                    16'h37FC: data_out = 8'hC5;
                    16'h37FD: data_out = 8'hC6;
                    16'h37FE: data_out = 8'hC7;
                    16'h37FF: data_out = 8'hC8;
                    16'h3800: data_out = 8'h38;
                    16'h3801: data_out = 8'h39;
                    16'h3802: data_out = 8'h3A;
                    16'h3803: data_out = 8'h3B;
                    16'h3804: data_out = 8'h3C;
                    16'h3805: data_out = 8'h3D;
                    16'h3806: data_out = 8'h3E;
                    16'h3807: data_out = 8'h3F;
                    16'h3808: data_out = 8'h40;
                    16'h3809: data_out = 8'h41;
                    16'h380A: data_out = 8'h42;
                    16'h380B: data_out = 8'h43;
                    16'h380C: data_out = 8'h44;
                    16'h380D: data_out = 8'h45;
                    16'h380E: data_out = 8'h46;
                    16'h380F: data_out = 8'h47;
                    16'h3810: data_out = 8'h48;
                    16'h3811: data_out = 8'h49;
                    16'h3812: data_out = 8'h4A;
                    16'h3813: data_out = 8'h4B;
                    16'h3814: data_out = 8'h4C;
                    16'h3815: data_out = 8'h4D;
                    16'h3816: data_out = 8'h4E;
                    16'h3817: data_out = 8'h4F;
                    16'h3818: data_out = 8'h50;
                    16'h3819: data_out = 8'h51;
                    16'h381A: data_out = 8'h52;
                    16'h381B: data_out = 8'h53;
                    16'h381C: data_out = 8'h54;
                    16'h381D: data_out = 8'h55;
                    16'h381E: data_out = 8'h56;
                    16'h381F: data_out = 8'h57;
                    16'h3820: data_out = 8'h58;
                    16'h3821: data_out = 8'h59;
                    16'h3822: data_out = 8'h5A;
                    16'h3823: data_out = 8'h5B;
                    16'h3824: data_out = 8'h5C;
                    16'h3825: data_out = 8'h5D;
                    16'h3826: data_out = 8'h5E;
                    16'h3827: data_out = 8'h5F;
                    16'h3828: data_out = 8'h60;
                    16'h3829: data_out = 8'h61;
                    16'h382A: data_out = 8'h62;
                    16'h382B: data_out = 8'h63;
                    16'h382C: data_out = 8'h64;
                    16'h382D: data_out = 8'h65;
                    16'h382E: data_out = 8'h66;
                    16'h382F: data_out = 8'h67;
                    16'h3830: data_out = 8'h68;
                    16'h3831: data_out = 8'h69;
                    16'h3832: data_out = 8'h6A;
                    16'h3833: data_out = 8'h6B;
                    16'h3834: data_out = 8'h6C;
                    16'h3835: data_out = 8'h6D;
                    16'h3836: data_out = 8'h6E;
                    16'h3837: data_out = 8'h6F;
                    16'h3838: data_out = 8'h70;
                    16'h3839: data_out = 8'h71;
                    16'h383A: data_out = 8'h72;
                    16'h383B: data_out = 8'h73;
                    16'h383C: data_out = 8'h74;
                    16'h383D: data_out = 8'h75;
                    16'h383E: data_out = 8'h76;
                    16'h383F: data_out = 8'h77;
                    16'h3840: data_out = 8'h78;
                    16'h3841: data_out = 8'h79;
                    16'h3842: data_out = 8'h7A;
                    16'h3843: data_out = 8'h7B;
                    16'h3844: data_out = 8'h7C;
                    16'h3845: data_out = 8'h7D;
                    16'h3846: data_out = 8'h7E;
                    16'h3847: data_out = 8'h7F;
                    16'h3848: data_out = 8'h80;
                    16'h3849: data_out = 8'h81;
                    16'h384A: data_out = 8'h82;
                    16'h384B: data_out = 8'h83;
                    16'h384C: data_out = 8'h84;
                    16'h384D: data_out = 8'h85;
                    16'h384E: data_out = 8'h86;
                    16'h384F: data_out = 8'h87;
                    16'h3850: data_out = 8'h88;
                    16'h3851: data_out = 8'h89;
                    16'h3852: data_out = 8'h8A;
                    16'h3853: data_out = 8'h8B;
                    16'h3854: data_out = 8'h8C;
                    16'h3855: data_out = 8'h8D;
                    16'h3856: data_out = 8'h8E;
                    16'h3857: data_out = 8'h8F;
                    16'h3858: data_out = 8'h90;
                    16'h3859: data_out = 8'h91;
                    16'h385A: data_out = 8'h92;
                    16'h385B: data_out = 8'h93;
                    16'h385C: data_out = 8'h94;
                    16'h385D: data_out = 8'h95;
                    16'h385E: data_out = 8'h96;
                    16'h385F: data_out = 8'h97;
                    16'h3860: data_out = 8'h98;
                    16'h3861: data_out = 8'h99;
                    16'h3862: data_out = 8'h9A;
                    16'h3863: data_out = 8'h9B;
                    16'h3864: data_out = 8'h9C;
                    16'h3865: data_out = 8'h9D;
                    16'h3866: data_out = 8'h9E;
                    16'h3867: data_out = 8'h9F;
                    16'h3868: data_out = 8'hA0;
                    16'h3869: data_out = 8'hA1;
                    16'h386A: data_out = 8'hA2;
                    16'h386B: data_out = 8'hA3;
                    16'h386C: data_out = 8'hA4;
                    16'h386D: data_out = 8'hA5;
                    16'h386E: data_out = 8'hA6;
                    16'h386F: data_out = 8'hA7;
                    16'h3870: data_out = 8'hA8;
                    16'h3871: data_out = 8'hA9;
                    16'h3872: data_out = 8'hAA;
                    16'h3873: data_out = 8'hAB;
                    16'h3874: data_out = 8'hAC;
                    16'h3875: data_out = 8'hAD;
                    16'h3876: data_out = 8'hAE;
                    16'h3877: data_out = 8'hAF;
                    16'h3878: data_out = 8'hB0;
                    16'h3879: data_out = 8'hB1;
                    16'h387A: data_out = 8'hB2;
                    16'h387B: data_out = 8'hB3;
                    16'h387C: data_out = 8'hB4;
                    16'h387D: data_out = 8'hB5;
                    16'h387E: data_out = 8'hB6;
                    16'h387F: data_out = 8'hB7;
                    16'h3880: data_out = 8'h38;
                    16'h3881: data_out = 8'h37;
                    16'h3882: data_out = 8'h36;
                    16'h3883: data_out = 8'h35;
                    16'h3884: data_out = 8'h34;
                    16'h3885: data_out = 8'h33;
                    16'h3886: data_out = 8'h32;
                    16'h3887: data_out = 8'h31;
                    16'h3888: data_out = 8'h30;
                    16'h3889: data_out = 8'h2F;
                    16'h388A: data_out = 8'h2E;
                    16'h388B: data_out = 8'h2D;
                    16'h388C: data_out = 8'h2C;
                    16'h388D: data_out = 8'h2B;
                    16'h388E: data_out = 8'h2A;
                    16'h388F: data_out = 8'h29;
                    16'h3890: data_out = 8'h28;
                    16'h3891: data_out = 8'h27;
                    16'h3892: data_out = 8'h26;
                    16'h3893: data_out = 8'h25;
                    16'h3894: data_out = 8'h24;
                    16'h3895: data_out = 8'h23;
                    16'h3896: data_out = 8'h22;
                    16'h3897: data_out = 8'h21;
                    16'h3898: data_out = 8'h20;
                    16'h3899: data_out = 8'h1F;
                    16'h389A: data_out = 8'h1E;
                    16'h389B: data_out = 8'h1D;
                    16'h389C: data_out = 8'h1C;
                    16'h389D: data_out = 8'h1B;
                    16'h389E: data_out = 8'h1A;
                    16'h389F: data_out = 8'h19;
                    16'h38A0: data_out = 8'h18;
                    16'h38A1: data_out = 8'h17;
                    16'h38A2: data_out = 8'h16;
                    16'h38A3: data_out = 8'h15;
                    16'h38A4: data_out = 8'h14;
                    16'h38A5: data_out = 8'h13;
                    16'h38A6: data_out = 8'h12;
                    16'h38A7: data_out = 8'h11;
                    16'h38A8: data_out = 8'h10;
                    16'h38A9: data_out = 8'hF;
                    16'h38AA: data_out = 8'hE;
                    16'h38AB: data_out = 8'hD;
                    16'h38AC: data_out = 8'hC;
                    16'h38AD: data_out = 8'hB;
                    16'h38AE: data_out = 8'hA;
                    16'h38AF: data_out = 8'h9;
                    16'h38B0: data_out = 8'h8;
                    16'h38B1: data_out = 8'h7;
                    16'h38B2: data_out = 8'h6;
                    16'h38B3: data_out = 8'h5;
                    16'h38B4: data_out = 8'h4;
                    16'h38B5: data_out = 8'h3;
                    16'h38B6: data_out = 8'h2;
                    16'h38B7: data_out = 8'h1;
                    16'h38B8: data_out = 8'h0;
                    16'h38B9: data_out = 8'h81;
                    16'h38BA: data_out = 8'h82;
                    16'h38BB: data_out = 8'h83;
                    16'h38BC: data_out = 8'h84;
                    16'h38BD: data_out = 8'h85;
                    16'h38BE: data_out = 8'h86;
                    16'h38BF: data_out = 8'h87;
                    16'h38C0: data_out = 8'h88;
                    16'h38C1: data_out = 8'h89;
                    16'h38C2: data_out = 8'h8A;
                    16'h38C3: data_out = 8'h8B;
                    16'h38C4: data_out = 8'h8C;
                    16'h38C5: data_out = 8'h8D;
                    16'h38C6: data_out = 8'h8E;
                    16'h38C7: data_out = 8'h8F;
                    16'h38C8: data_out = 8'h90;
                    16'h38C9: data_out = 8'h91;
                    16'h38CA: data_out = 8'h92;
                    16'h38CB: data_out = 8'h93;
                    16'h38CC: data_out = 8'h94;
                    16'h38CD: data_out = 8'h95;
                    16'h38CE: data_out = 8'h96;
                    16'h38CF: data_out = 8'h97;
                    16'h38D0: data_out = 8'h98;
                    16'h38D1: data_out = 8'h99;
                    16'h38D2: data_out = 8'h9A;
                    16'h38D3: data_out = 8'h9B;
                    16'h38D4: data_out = 8'h9C;
                    16'h38D5: data_out = 8'h9D;
                    16'h38D6: data_out = 8'h9E;
                    16'h38D7: data_out = 8'h9F;
                    16'h38D8: data_out = 8'hA0;
                    16'h38D9: data_out = 8'hA1;
                    16'h38DA: data_out = 8'hA2;
                    16'h38DB: data_out = 8'hA3;
                    16'h38DC: data_out = 8'hA4;
                    16'h38DD: data_out = 8'hA5;
                    16'h38DE: data_out = 8'hA6;
                    16'h38DF: data_out = 8'hA7;
                    16'h38E0: data_out = 8'hA8;
                    16'h38E1: data_out = 8'hA9;
                    16'h38E2: data_out = 8'hAA;
                    16'h38E3: data_out = 8'hAB;
                    16'h38E4: data_out = 8'hAC;
                    16'h38E5: data_out = 8'hAD;
                    16'h38E6: data_out = 8'hAE;
                    16'h38E7: data_out = 8'hAF;
                    16'h38E8: data_out = 8'hB0;
                    16'h38E9: data_out = 8'hB1;
                    16'h38EA: data_out = 8'hB2;
                    16'h38EB: data_out = 8'hB3;
                    16'h38EC: data_out = 8'hB4;
                    16'h38ED: data_out = 8'hB5;
                    16'h38EE: data_out = 8'hB6;
                    16'h38EF: data_out = 8'hB7;
                    16'h38F0: data_out = 8'hB8;
                    16'h38F1: data_out = 8'hB9;
                    16'h38F2: data_out = 8'hBA;
                    16'h38F3: data_out = 8'hBB;
                    16'h38F4: data_out = 8'hBC;
                    16'h38F5: data_out = 8'hBD;
                    16'h38F6: data_out = 8'hBE;
                    16'h38F7: data_out = 8'hBF;
                    16'h38F8: data_out = 8'hC0;
                    16'h38F9: data_out = 8'hC1;
                    16'h38FA: data_out = 8'hC2;
                    16'h38FB: data_out = 8'hC3;
                    16'h38FC: data_out = 8'hC4;
                    16'h38FD: data_out = 8'hC5;
                    16'h38FE: data_out = 8'hC6;
                    16'h38FF: data_out = 8'hC7;
                    16'h3900: data_out = 8'h39;
                    16'h3901: data_out = 8'h3A;
                    16'h3902: data_out = 8'h3B;
                    16'h3903: data_out = 8'h3C;
                    16'h3904: data_out = 8'h3D;
                    16'h3905: data_out = 8'h3E;
                    16'h3906: data_out = 8'h3F;
                    16'h3907: data_out = 8'h40;
                    16'h3908: data_out = 8'h41;
                    16'h3909: data_out = 8'h42;
                    16'h390A: data_out = 8'h43;
                    16'h390B: data_out = 8'h44;
                    16'h390C: data_out = 8'h45;
                    16'h390D: data_out = 8'h46;
                    16'h390E: data_out = 8'h47;
                    16'h390F: data_out = 8'h48;
                    16'h3910: data_out = 8'h49;
                    16'h3911: data_out = 8'h4A;
                    16'h3912: data_out = 8'h4B;
                    16'h3913: data_out = 8'h4C;
                    16'h3914: data_out = 8'h4D;
                    16'h3915: data_out = 8'h4E;
                    16'h3916: data_out = 8'h4F;
                    16'h3917: data_out = 8'h50;
                    16'h3918: data_out = 8'h51;
                    16'h3919: data_out = 8'h52;
                    16'h391A: data_out = 8'h53;
                    16'h391B: data_out = 8'h54;
                    16'h391C: data_out = 8'h55;
                    16'h391D: data_out = 8'h56;
                    16'h391E: data_out = 8'h57;
                    16'h391F: data_out = 8'h58;
                    16'h3920: data_out = 8'h59;
                    16'h3921: data_out = 8'h5A;
                    16'h3922: data_out = 8'h5B;
                    16'h3923: data_out = 8'h5C;
                    16'h3924: data_out = 8'h5D;
                    16'h3925: data_out = 8'h5E;
                    16'h3926: data_out = 8'h5F;
                    16'h3927: data_out = 8'h60;
                    16'h3928: data_out = 8'h61;
                    16'h3929: data_out = 8'h62;
                    16'h392A: data_out = 8'h63;
                    16'h392B: data_out = 8'h64;
                    16'h392C: data_out = 8'h65;
                    16'h392D: data_out = 8'h66;
                    16'h392E: data_out = 8'h67;
                    16'h392F: data_out = 8'h68;
                    16'h3930: data_out = 8'h69;
                    16'h3931: data_out = 8'h6A;
                    16'h3932: data_out = 8'h6B;
                    16'h3933: data_out = 8'h6C;
                    16'h3934: data_out = 8'h6D;
                    16'h3935: data_out = 8'h6E;
                    16'h3936: data_out = 8'h6F;
                    16'h3937: data_out = 8'h70;
                    16'h3938: data_out = 8'h71;
                    16'h3939: data_out = 8'h72;
                    16'h393A: data_out = 8'h73;
                    16'h393B: data_out = 8'h74;
                    16'h393C: data_out = 8'h75;
                    16'h393D: data_out = 8'h76;
                    16'h393E: data_out = 8'h77;
                    16'h393F: data_out = 8'h78;
                    16'h3940: data_out = 8'h79;
                    16'h3941: data_out = 8'h7A;
                    16'h3942: data_out = 8'h7B;
                    16'h3943: data_out = 8'h7C;
                    16'h3944: data_out = 8'h7D;
                    16'h3945: data_out = 8'h7E;
                    16'h3946: data_out = 8'h7F;
                    16'h3947: data_out = 8'h80;
                    16'h3948: data_out = 8'h81;
                    16'h3949: data_out = 8'h82;
                    16'h394A: data_out = 8'h83;
                    16'h394B: data_out = 8'h84;
                    16'h394C: data_out = 8'h85;
                    16'h394D: data_out = 8'h86;
                    16'h394E: data_out = 8'h87;
                    16'h394F: data_out = 8'h88;
                    16'h3950: data_out = 8'h89;
                    16'h3951: data_out = 8'h8A;
                    16'h3952: data_out = 8'h8B;
                    16'h3953: data_out = 8'h8C;
                    16'h3954: data_out = 8'h8D;
                    16'h3955: data_out = 8'h8E;
                    16'h3956: data_out = 8'h8F;
                    16'h3957: data_out = 8'h90;
                    16'h3958: data_out = 8'h91;
                    16'h3959: data_out = 8'h92;
                    16'h395A: data_out = 8'h93;
                    16'h395B: data_out = 8'h94;
                    16'h395C: data_out = 8'h95;
                    16'h395D: data_out = 8'h96;
                    16'h395E: data_out = 8'h97;
                    16'h395F: data_out = 8'h98;
                    16'h3960: data_out = 8'h99;
                    16'h3961: data_out = 8'h9A;
                    16'h3962: data_out = 8'h9B;
                    16'h3963: data_out = 8'h9C;
                    16'h3964: data_out = 8'h9D;
                    16'h3965: data_out = 8'h9E;
                    16'h3966: data_out = 8'h9F;
                    16'h3967: data_out = 8'hA0;
                    16'h3968: data_out = 8'hA1;
                    16'h3969: data_out = 8'hA2;
                    16'h396A: data_out = 8'hA3;
                    16'h396B: data_out = 8'hA4;
                    16'h396C: data_out = 8'hA5;
                    16'h396D: data_out = 8'hA6;
                    16'h396E: data_out = 8'hA7;
                    16'h396F: data_out = 8'hA8;
                    16'h3970: data_out = 8'hA9;
                    16'h3971: data_out = 8'hAA;
                    16'h3972: data_out = 8'hAB;
                    16'h3973: data_out = 8'hAC;
                    16'h3974: data_out = 8'hAD;
                    16'h3975: data_out = 8'hAE;
                    16'h3976: data_out = 8'hAF;
                    16'h3977: data_out = 8'hB0;
                    16'h3978: data_out = 8'hB1;
                    16'h3979: data_out = 8'hB2;
                    16'h397A: data_out = 8'hB3;
                    16'h397B: data_out = 8'hB4;
                    16'h397C: data_out = 8'hB5;
                    16'h397D: data_out = 8'hB6;
                    16'h397E: data_out = 8'hB7;
                    16'h397F: data_out = 8'hB8;
                    16'h3980: data_out = 8'h39;
                    16'h3981: data_out = 8'h38;
                    16'h3982: data_out = 8'h37;
                    16'h3983: data_out = 8'h36;
                    16'h3984: data_out = 8'h35;
                    16'h3985: data_out = 8'h34;
                    16'h3986: data_out = 8'h33;
                    16'h3987: data_out = 8'h32;
                    16'h3988: data_out = 8'h31;
                    16'h3989: data_out = 8'h30;
                    16'h398A: data_out = 8'h2F;
                    16'h398B: data_out = 8'h2E;
                    16'h398C: data_out = 8'h2D;
                    16'h398D: data_out = 8'h2C;
                    16'h398E: data_out = 8'h2B;
                    16'h398F: data_out = 8'h2A;
                    16'h3990: data_out = 8'h29;
                    16'h3991: data_out = 8'h28;
                    16'h3992: data_out = 8'h27;
                    16'h3993: data_out = 8'h26;
                    16'h3994: data_out = 8'h25;
                    16'h3995: data_out = 8'h24;
                    16'h3996: data_out = 8'h23;
                    16'h3997: data_out = 8'h22;
                    16'h3998: data_out = 8'h21;
                    16'h3999: data_out = 8'h20;
                    16'h399A: data_out = 8'h1F;
                    16'h399B: data_out = 8'h1E;
                    16'h399C: data_out = 8'h1D;
                    16'h399D: data_out = 8'h1C;
                    16'h399E: data_out = 8'h1B;
                    16'h399F: data_out = 8'h1A;
                    16'h39A0: data_out = 8'h19;
                    16'h39A1: data_out = 8'h18;
                    16'h39A2: data_out = 8'h17;
                    16'h39A3: data_out = 8'h16;
                    16'h39A4: data_out = 8'h15;
                    16'h39A5: data_out = 8'h14;
                    16'h39A6: data_out = 8'h13;
                    16'h39A7: data_out = 8'h12;
                    16'h39A8: data_out = 8'h11;
                    16'h39A9: data_out = 8'h10;
                    16'h39AA: data_out = 8'hF;
                    16'h39AB: data_out = 8'hE;
                    16'h39AC: data_out = 8'hD;
                    16'h39AD: data_out = 8'hC;
                    16'h39AE: data_out = 8'hB;
                    16'h39AF: data_out = 8'hA;
                    16'h39B0: data_out = 8'h9;
                    16'h39B1: data_out = 8'h8;
                    16'h39B2: data_out = 8'h7;
                    16'h39B3: data_out = 8'h6;
                    16'h39B4: data_out = 8'h5;
                    16'h39B5: data_out = 8'h4;
                    16'h39B6: data_out = 8'h3;
                    16'h39B7: data_out = 8'h2;
                    16'h39B8: data_out = 8'h1;
                    16'h39B9: data_out = 8'h0;
                    16'h39BA: data_out = 8'h81;
                    16'h39BB: data_out = 8'h82;
                    16'h39BC: data_out = 8'h83;
                    16'h39BD: data_out = 8'h84;
                    16'h39BE: data_out = 8'h85;
                    16'h39BF: data_out = 8'h86;
                    16'h39C0: data_out = 8'h87;
                    16'h39C1: data_out = 8'h88;
                    16'h39C2: data_out = 8'h89;
                    16'h39C3: data_out = 8'h8A;
                    16'h39C4: data_out = 8'h8B;
                    16'h39C5: data_out = 8'h8C;
                    16'h39C6: data_out = 8'h8D;
                    16'h39C7: data_out = 8'h8E;
                    16'h39C8: data_out = 8'h8F;
                    16'h39C9: data_out = 8'h90;
                    16'h39CA: data_out = 8'h91;
                    16'h39CB: data_out = 8'h92;
                    16'h39CC: data_out = 8'h93;
                    16'h39CD: data_out = 8'h94;
                    16'h39CE: data_out = 8'h95;
                    16'h39CF: data_out = 8'h96;
                    16'h39D0: data_out = 8'h97;
                    16'h39D1: data_out = 8'h98;
                    16'h39D2: data_out = 8'h99;
                    16'h39D3: data_out = 8'h9A;
                    16'h39D4: data_out = 8'h9B;
                    16'h39D5: data_out = 8'h9C;
                    16'h39D6: data_out = 8'h9D;
                    16'h39D7: data_out = 8'h9E;
                    16'h39D8: data_out = 8'h9F;
                    16'h39D9: data_out = 8'hA0;
                    16'h39DA: data_out = 8'hA1;
                    16'h39DB: data_out = 8'hA2;
                    16'h39DC: data_out = 8'hA3;
                    16'h39DD: data_out = 8'hA4;
                    16'h39DE: data_out = 8'hA5;
                    16'h39DF: data_out = 8'hA6;
                    16'h39E0: data_out = 8'hA7;
                    16'h39E1: data_out = 8'hA8;
                    16'h39E2: data_out = 8'hA9;
                    16'h39E3: data_out = 8'hAA;
                    16'h39E4: data_out = 8'hAB;
                    16'h39E5: data_out = 8'hAC;
                    16'h39E6: data_out = 8'hAD;
                    16'h39E7: data_out = 8'hAE;
                    16'h39E8: data_out = 8'hAF;
                    16'h39E9: data_out = 8'hB0;
                    16'h39EA: data_out = 8'hB1;
                    16'h39EB: data_out = 8'hB2;
                    16'h39EC: data_out = 8'hB3;
                    16'h39ED: data_out = 8'hB4;
                    16'h39EE: data_out = 8'hB5;
                    16'h39EF: data_out = 8'hB6;
                    16'h39F0: data_out = 8'hB7;
                    16'h39F1: data_out = 8'hB8;
                    16'h39F2: data_out = 8'hB9;
                    16'h39F3: data_out = 8'hBA;
                    16'h39F4: data_out = 8'hBB;
                    16'h39F5: data_out = 8'hBC;
                    16'h39F6: data_out = 8'hBD;
                    16'h39F7: data_out = 8'hBE;
                    16'h39F8: data_out = 8'hBF;
                    16'h39F9: data_out = 8'hC0;
                    16'h39FA: data_out = 8'hC1;
                    16'h39FB: data_out = 8'hC2;
                    16'h39FC: data_out = 8'hC3;
                    16'h39FD: data_out = 8'hC4;
                    16'h39FE: data_out = 8'hC5;
                    16'h39FF: data_out = 8'hC6;
                    16'h3A00: data_out = 8'h3A;
                    16'h3A01: data_out = 8'h3B;
                    16'h3A02: data_out = 8'h3C;
                    16'h3A03: data_out = 8'h3D;
                    16'h3A04: data_out = 8'h3E;
                    16'h3A05: data_out = 8'h3F;
                    16'h3A06: data_out = 8'h40;
                    16'h3A07: data_out = 8'h41;
                    16'h3A08: data_out = 8'h42;
                    16'h3A09: data_out = 8'h43;
                    16'h3A0A: data_out = 8'h44;
                    16'h3A0B: data_out = 8'h45;
                    16'h3A0C: data_out = 8'h46;
                    16'h3A0D: data_out = 8'h47;
                    16'h3A0E: data_out = 8'h48;
                    16'h3A0F: data_out = 8'h49;
                    16'h3A10: data_out = 8'h4A;
                    16'h3A11: data_out = 8'h4B;
                    16'h3A12: data_out = 8'h4C;
                    16'h3A13: data_out = 8'h4D;
                    16'h3A14: data_out = 8'h4E;
                    16'h3A15: data_out = 8'h4F;
                    16'h3A16: data_out = 8'h50;
                    16'h3A17: data_out = 8'h51;
                    16'h3A18: data_out = 8'h52;
                    16'h3A19: data_out = 8'h53;
                    16'h3A1A: data_out = 8'h54;
                    16'h3A1B: data_out = 8'h55;
                    16'h3A1C: data_out = 8'h56;
                    16'h3A1D: data_out = 8'h57;
                    16'h3A1E: data_out = 8'h58;
                    16'h3A1F: data_out = 8'h59;
                    16'h3A20: data_out = 8'h5A;
                    16'h3A21: data_out = 8'h5B;
                    16'h3A22: data_out = 8'h5C;
                    16'h3A23: data_out = 8'h5D;
                    16'h3A24: data_out = 8'h5E;
                    16'h3A25: data_out = 8'h5F;
                    16'h3A26: data_out = 8'h60;
                    16'h3A27: data_out = 8'h61;
                    16'h3A28: data_out = 8'h62;
                    16'h3A29: data_out = 8'h63;
                    16'h3A2A: data_out = 8'h64;
                    16'h3A2B: data_out = 8'h65;
                    16'h3A2C: data_out = 8'h66;
                    16'h3A2D: data_out = 8'h67;
                    16'h3A2E: data_out = 8'h68;
                    16'h3A2F: data_out = 8'h69;
                    16'h3A30: data_out = 8'h6A;
                    16'h3A31: data_out = 8'h6B;
                    16'h3A32: data_out = 8'h6C;
                    16'h3A33: data_out = 8'h6D;
                    16'h3A34: data_out = 8'h6E;
                    16'h3A35: data_out = 8'h6F;
                    16'h3A36: data_out = 8'h70;
                    16'h3A37: data_out = 8'h71;
                    16'h3A38: data_out = 8'h72;
                    16'h3A39: data_out = 8'h73;
                    16'h3A3A: data_out = 8'h74;
                    16'h3A3B: data_out = 8'h75;
                    16'h3A3C: data_out = 8'h76;
                    16'h3A3D: data_out = 8'h77;
                    16'h3A3E: data_out = 8'h78;
                    16'h3A3F: data_out = 8'h79;
                    16'h3A40: data_out = 8'h7A;
                    16'h3A41: data_out = 8'h7B;
                    16'h3A42: data_out = 8'h7C;
                    16'h3A43: data_out = 8'h7D;
                    16'h3A44: data_out = 8'h7E;
                    16'h3A45: data_out = 8'h7F;
                    16'h3A46: data_out = 8'h80;
                    16'h3A47: data_out = 8'h81;
                    16'h3A48: data_out = 8'h82;
                    16'h3A49: data_out = 8'h83;
                    16'h3A4A: data_out = 8'h84;
                    16'h3A4B: data_out = 8'h85;
                    16'h3A4C: data_out = 8'h86;
                    16'h3A4D: data_out = 8'h87;
                    16'h3A4E: data_out = 8'h88;
                    16'h3A4F: data_out = 8'h89;
                    16'h3A50: data_out = 8'h8A;
                    16'h3A51: data_out = 8'h8B;
                    16'h3A52: data_out = 8'h8C;
                    16'h3A53: data_out = 8'h8D;
                    16'h3A54: data_out = 8'h8E;
                    16'h3A55: data_out = 8'h8F;
                    16'h3A56: data_out = 8'h90;
                    16'h3A57: data_out = 8'h91;
                    16'h3A58: data_out = 8'h92;
                    16'h3A59: data_out = 8'h93;
                    16'h3A5A: data_out = 8'h94;
                    16'h3A5B: data_out = 8'h95;
                    16'h3A5C: data_out = 8'h96;
                    16'h3A5D: data_out = 8'h97;
                    16'h3A5E: data_out = 8'h98;
                    16'h3A5F: data_out = 8'h99;
                    16'h3A60: data_out = 8'h9A;
                    16'h3A61: data_out = 8'h9B;
                    16'h3A62: data_out = 8'h9C;
                    16'h3A63: data_out = 8'h9D;
                    16'h3A64: data_out = 8'h9E;
                    16'h3A65: data_out = 8'h9F;
                    16'h3A66: data_out = 8'hA0;
                    16'h3A67: data_out = 8'hA1;
                    16'h3A68: data_out = 8'hA2;
                    16'h3A69: data_out = 8'hA3;
                    16'h3A6A: data_out = 8'hA4;
                    16'h3A6B: data_out = 8'hA5;
                    16'h3A6C: data_out = 8'hA6;
                    16'h3A6D: data_out = 8'hA7;
                    16'h3A6E: data_out = 8'hA8;
                    16'h3A6F: data_out = 8'hA9;
                    16'h3A70: data_out = 8'hAA;
                    16'h3A71: data_out = 8'hAB;
                    16'h3A72: data_out = 8'hAC;
                    16'h3A73: data_out = 8'hAD;
                    16'h3A74: data_out = 8'hAE;
                    16'h3A75: data_out = 8'hAF;
                    16'h3A76: data_out = 8'hB0;
                    16'h3A77: data_out = 8'hB1;
                    16'h3A78: data_out = 8'hB2;
                    16'h3A79: data_out = 8'hB3;
                    16'h3A7A: data_out = 8'hB4;
                    16'h3A7B: data_out = 8'hB5;
                    16'h3A7C: data_out = 8'hB6;
                    16'h3A7D: data_out = 8'hB7;
                    16'h3A7E: data_out = 8'hB8;
                    16'h3A7F: data_out = 8'hB9;
                    16'h3A80: data_out = 8'h3A;
                    16'h3A81: data_out = 8'h39;
                    16'h3A82: data_out = 8'h38;
                    16'h3A83: data_out = 8'h37;
                    16'h3A84: data_out = 8'h36;
                    16'h3A85: data_out = 8'h35;
                    16'h3A86: data_out = 8'h34;
                    16'h3A87: data_out = 8'h33;
                    16'h3A88: data_out = 8'h32;
                    16'h3A89: data_out = 8'h31;
                    16'h3A8A: data_out = 8'h30;
                    16'h3A8B: data_out = 8'h2F;
                    16'h3A8C: data_out = 8'h2E;
                    16'h3A8D: data_out = 8'h2D;
                    16'h3A8E: data_out = 8'h2C;
                    16'h3A8F: data_out = 8'h2B;
                    16'h3A90: data_out = 8'h2A;
                    16'h3A91: data_out = 8'h29;
                    16'h3A92: data_out = 8'h28;
                    16'h3A93: data_out = 8'h27;
                    16'h3A94: data_out = 8'h26;
                    16'h3A95: data_out = 8'h25;
                    16'h3A96: data_out = 8'h24;
                    16'h3A97: data_out = 8'h23;
                    16'h3A98: data_out = 8'h22;
                    16'h3A99: data_out = 8'h21;
                    16'h3A9A: data_out = 8'h20;
                    16'h3A9B: data_out = 8'h1F;
                    16'h3A9C: data_out = 8'h1E;
                    16'h3A9D: data_out = 8'h1D;
                    16'h3A9E: data_out = 8'h1C;
                    16'h3A9F: data_out = 8'h1B;
                    16'h3AA0: data_out = 8'h1A;
                    16'h3AA1: data_out = 8'h19;
                    16'h3AA2: data_out = 8'h18;
                    16'h3AA3: data_out = 8'h17;
                    16'h3AA4: data_out = 8'h16;
                    16'h3AA5: data_out = 8'h15;
                    16'h3AA6: data_out = 8'h14;
                    16'h3AA7: data_out = 8'h13;
                    16'h3AA8: data_out = 8'h12;
                    16'h3AA9: data_out = 8'h11;
                    16'h3AAA: data_out = 8'h10;
                    16'h3AAB: data_out = 8'hF;
                    16'h3AAC: data_out = 8'hE;
                    16'h3AAD: data_out = 8'hD;
                    16'h3AAE: data_out = 8'hC;
                    16'h3AAF: data_out = 8'hB;
                    16'h3AB0: data_out = 8'hA;
                    16'h3AB1: data_out = 8'h9;
                    16'h3AB2: data_out = 8'h8;
                    16'h3AB3: data_out = 8'h7;
                    16'h3AB4: data_out = 8'h6;
                    16'h3AB5: data_out = 8'h5;
                    16'h3AB6: data_out = 8'h4;
                    16'h3AB7: data_out = 8'h3;
                    16'h3AB8: data_out = 8'h2;
                    16'h3AB9: data_out = 8'h1;
                    16'h3ABA: data_out = 8'h0;
                    16'h3ABB: data_out = 8'h81;
                    16'h3ABC: data_out = 8'h82;
                    16'h3ABD: data_out = 8'h83;
                    16'h3ABE: data_out = 8'h84;
                    16'h3ABF: data_out = 8'h85;
                    16'h3AC0: data_out = 8'h86;
                    16'h3AC1: data_out = 8'h87;
                    16'h3AC2: data_out = 8'h88;
                    16'h3AC3: data_out = 8'h89;
                    16'h3AC4: data_out = 8'h8A;
                    16'h3AC5: data_out = 8'h8B;
                    16'h3AC6: data_out = 8'h8C;
                    16'h3AC7: data_out = 8'h8D;
                    16'h3AC8: data_out = 8'h8E;
                    16'h3AC9: data_out = 8'h8F;
                    16'h3ACA: data_out = 8'h90;
                    16'h3ACB: data_out = 8'h91;
                    16'h3ACC: data_out = 8'h92;
                    16'h3ACD: data_out = 8'h93;
                    16'h3ACE: data_out = 8'h94;
                    16'h3ACF: data_out = 8'h95;
                    16'h3AD0: data_out = 8'h96;
                    16'h3AD1: data_out = 8'h97;
                    16'h3AD2: data_out = 8'h98;
                    16'h3AD3: data_out = 8'h99;
                    16'h3AD4: data_out = 8'h9A;
                    16'h3AD5: data_out = 8'h9B;
                    16'h3AD6: data_out = 8'h9C;
                    16'h3AD7: data_out = 8'h9D;
                    16'h3AD8: data_out = 8'h9E;
                    16'h3AD9: data_out = 8'h9F;
                    16'h3ADA: data_out = 8'hA0;
                    16'h3ADB: data_out = 8'hA1;
                    16'h3ADC: data_out = 8'hA2;
                    16'h3ADD: data_out = 8'hA3;
                    16'h3ADE: data_out = 8'hA4;
                    16'h3ADF: data_out = 8'hA5;
                    16'h3AE0: data_out = 8'hA6;
                    16'h3AE1: data_out = 8'hA7;
                    16'h3AE2: data_out = 8'hA8;
                    16'h3AE3: data_out = 8'hA9;
                    16'h3AE4: data_out = 8'hAA;
                    16'h3AE5: data_out = 8'hAB;
                    16'h3AE6: data_out = 8'hAC;
                    16'h3AE7: data_out = 8'hAD;
                    16'h3AE8: data_out = 8'hAE;
                    16'h3AE9: data_out = 8'hAF;
                    16'h3AEA: data_out = 8'hB0;
                    16'h3AEB: data_out = 8'hB1;
                    16'h3AEC: data_out = 8'hB2;
                    16'h3AED: data_out = 8'hB3;
                    16'h3AEE: data_out = 8'hB4;
                    16'h3AEF: data_out = 8'hB5;
                    16'h3AF0: data_out = 8'hB6;
                    16'h3AF1: data_out = 8'hB7;
                    16'h3AF2: data_out = 8'hB8;
                    16'h3AF3: data_out = 8'hB9;
                    16'h3AF4: data_out = 8'hBA;
                    16'h3AF5: data_out = 8'hBB;
                    16'h3AF6: data_out = 8'hBC;
                    16'h3AF7: data_out = 8'hBD;
                    16'h3AF8: data_out = 8'hBE;
                    16'h3AF9: data_out = 8'hBF;
                    16'h3AFA: data_out = 8'hC0;
                    16'h3AFB: data_out = 8'hC1;
                    16'h3AFC: data_out = 8'hC2;
                    16'h3AFD: data_out = 8'hC3;
                    16'h3AFE: data_out = 8'hC4;
                    16'h3AFF: data_out = 8'hC5;
                    16'h3B00: data_out = 8'h3B;
                    16'h3B01: data_out = 8'h3C;
                    16'h3B02: data_out = 8'h3D;
                    16'h3B03: data_out = 8'h3E;
                    16'h3B04: data_out = 8'h3F;
                    16'h3B05: data_out = 8'h40;
                    16'h3B06: data_out = 8'h41;
                    16'h3B07: data_out = 8'h42;
                    16'h3B08: data_out = 8'h43;
                    16'h3B09: data_out = 8'h44;
                    16'h3B0A: data_out = 8'h45;
                    16'h3B0B: data_out = 8'h46;
                    16'h3B0C: data_out = 8'h47;
                    16'h3B0D: data_out = 8'h48;
                    16'h3B0E: data_out = 8'h49;
                    16'h3B0F: data_out = 8'h4A;
                    16'h3B10: data_out = 8'h4B;
                    16'h3B11: data_out = 8'h4C;
                    16'h3B12: data_out = 8'h4D;
                    16'h3B13: data_out = 8'h4E;
                    16'h3B14: data_out = 8'h4F;
                    16'h3B15: data_out = 8'h50;
                    16'h3B16: data_out = 8'h51;
                    16'h3B17: data_out = 8'h52;
                    16'h3B18: data_out = 8'h53;
                    16'h3B19: data_out = 8'h54;
                    16'h3B1A: data_out = 8'h55;
                    16'h3B1B: data_out = 8'h56;
                    16'h3B1C: data_out = 8'h57;
                    16'h3B1D: data_out = 8'h58;
                    16'h3B1E: data_out = 8'h59;
                    16'h3B1F: data_out = 8'h5A;
                    16'h3B20: data_out = 8'h5B;
                    16'h3B21: data_out = 8'h5C;
                    16'h3B22: data_out = 8'h5D;
                    16'h3B23: data_out = 8'h5E;
                    16'h3B24: data_out = 8'h5F;
                    16'h3B25: data_out = 8'h60;
                    16'h3B26: data_out = 8'h61;
                    16'h3B27: data_out = 8'h62;
                    16'h3B28: data_out = 8'h63;
                    16'h3B29: data_out = 8'h64;
                    16'h3B2A: data_out = 8'h65;
                    16'h3B2B: data_out = 8'h66;
                    16'h3B2C: data_out = 8'h67;
                    16'h3B2D: data_out = 8'h68;
                    16'h3B2E: data_out = 8'h69;
                    16'h3B2F: data_out = 8'h6A;
                    16'h3B30: data_out = 8'h6B;
                    16'h3B31: data_out = 8'h6C;
                    16'h3B32: data_out = 8'h6D;
                    16'h3B33: data_out = 8'h6E;
                    16'h3B34: data_out = 8'h6F;
                    16'h3B35: data_out = 8'h70;
                    16'h3B36: data_out = 8'h71;
                    16'h3B37: data_out = 8'h72;
                    16'h3B38: data_out = 8'h73;
                    16'h3B39: data_out = 8'h74;
                    16'h3B3A: data_out = 8'h75;
                    16'h3B3B: data_out = 8'h76;
                    16'h3B3C: data_out = 8'h77;
                    16'h3B3D: data_out = 8'h78;
                    16'h3B3E: data_out = 8'h79;
                    16'h3B3F: data_out = 8'h7A;
                    16'h3B40: data_out = 8'h7B;
                    16'h3B41: data_out = 8'h7C;
                    16'h3B42: data_out = 8'h7D;
                    16'h3B43: data_out = 8'h7E;
                    16'h3B44: data_out = 8'h7F;
                    16'h3B45: data_out = 8'h80;
                    16'h3B46: data_out = 8'h81;
                    16'h3B47: data_out = 8'h82;
                    16'h3B48: data_out = 8'h83;
                    16'h3B49: data_out = 8'h84;
                    16'h3B4A: data_out = 8'h85;
                    16'h3B4B: data_out = 8'h86;
                    16'h3B4C: data_out = 8'h87;
                    16'h3B4D: data_out = 8'h88;
                    16'h3B4E: data_out = 8'h89;
                    16'h3B4F: data_out = 8'h8A;
                    16'h3B50: data_out = 8'h8B;
                    16'h3B51: data_out = 8'h8C;
                    16'h3B52: data_out = 8'h8D;
                    16'h3B53: data_out = 8'h8E;
                    16'h3B54: data_out = 8'h8F;
                    16'h3B55: data_out = 8'h90;
                    16'h3B56: data_out = 8'h91;
                    16'h3B57: data_out = 8'h92;
                    16'h3B58: data_out = 8'h93;
                    16'h3B59: data_out = 8'h94;
                    16'h3B5A: data_out = 8'h95;
                    16'h3B5B: data_out = 8'h96;
                    16'h3B5C: data_out = 8'h97;
                    16'h3B5D: data_out = 8'h98;
                    16'h3B5E: data_out = 8'h99;
                    16'h3B5F: data_out = 8'h9A;
                    16'h3B60: data_out = 8'h9B;
                    16'h3B61: data_out = 8'h9C;
                    16'h3B62: data_out = 8'h9D;
                    16'h3B63: data_out = 8'h9E;
                    16'h3B64: data_out = 8'h9F;
                    16'h3B65: data_out = 8'hA0;
                    16'h3B66: data_out = 8'hA1;
                    16'h3B67: data_out = 8'hA2;
                    16'h3B68: data_out = 8'hA3;
                    16'h3B69: data_out = 8'hA4;
                    16'h3B6A: data_out = 8'hA5;
                    16'h3B6B: data_out = 8'hA6;
                    16'h3B6C: data_out = 8'hA7;
                    16'h3B6D: data_out = 8'hA8;
                    16'h3B6E: data_out = 8'hA9;
                    16'h3B6F: data_out = 8'hAA;
                    16'h3B70: data_out = 8'hAB;
                    16'h3B71: data_out = 8'hAC;
                    16'h3B72: data_out = 8'hAD;
                    16'h3B73: data_out = 8'hAE;
                    16'h3B74: data_out = 8'hAF;
                    16'h3B75: data_out = 8'hB0;
                    16'h3B76: data_out = 8'hB1;
                    16'h3B77: data_out = 8'hB2;
                    16'h3B78: data_out = 8'hB3;
                    16'h3B79: data_out = 8'hB4;
                    16'h3B7A: data_out = 8'hB5;
                    16'h3B7B: data_out = 8'hB6;
                    16'h3B7C: data_out = 8'hB7;
                    16'h3B7D: data_out = 8'hB8;
                    16'h3B7E: data_out = 8'hB9;
                    16'h3B7F: data_out = 8'hBA;
                    16'h3B80: data_out = 8'h3B;
                    16'h3B81: data_out = 8'h3A;
                    16'h3B82: data_out = 8'h39;
                    16'h3B83: data_out = 8'h38;
                    16'h3B84: data_out = 8'h37;
                    16'h3B85: data_out = 8'h36;
                    16'h3B86: data_out = 8'h35;
                    16'h3B87: data_out = 8'h34;
                    16'h3B88: data_out = 8'h33;
                    16'h3B89: data_out = 8'h32;
                    16'h3B8A: data_out = 8'h31;
                    16'h3B8B: data_out = 8'h30;
                    16'h3B8C: data_out = 8'h2F;
                    16'h3B8D: data_out = 8'h2E;
                    16'h3B8E: data_out = 8'h2D;
                    16'h3B8F: data_out = 8'h2C;
                    16'h3B90: data_out = 8'h2B;
                    16'h3B91: data_out = 8'h2A;
                    16'h3B92: data_out = 8'h29;
                    16'h3B93: data_out = 8'h28;
                    16'h3B94: data_out = 8'h27;
                    16'h3B95: data_out = 8'h26;
                    16'h3B96: data_out = 8'h25;
                    16'h3B97: data_out = 8'h24;
                    16'h3B98: data_out = 8'h23;
                    16'h3B99: data_out = 8'h22;
                    16'h3B9A: data_out = 8'h21;
                    16'h3B9B: data_out = 8'h20;
                    16'h3B9C: data_out = 8'h1F;
                    16'h3B9D: data_out = 8'h1E;
                    16'h3B9E: data_out = 8'h1D;
                    16'h3B9F: data_out = 8'h1C;
                    16'h3BA0: data_out = 8'h1B;
                    16'h3BA1: data_out = 8'h1A;
                    16'h3BA2: data_out = 8'h19;
                    16'h3BA3: data_out = 8'h18;
                    16'h3BA4: data_out = 8'h17;
                    16'h3BA5: data_out = 8'h16;
                    16'h3BA6: data_out = 8'h15;
                    16'h3BA7: data_out = 8'h14;
                    16'h3BA8: data_out = 8'h13;
                    16'h3BA9: data_out = 8'h12;
                    16'h3BAA: data_out = 8'h11;
                    16'h3BAB: data_out = 8'h10;
                    16'h3BAC: data_out = 8'hF;
                    16'h3BAD: data_out = 8'hE;
                    16'h3BAE: data_out = 8'hD;
                    16'h3BAF: data_out = 8'hC;
                    16'h3BB0: data_out = 8'hB;
                    16'h3BB1: data_out = 8'hA;
                    16'h3BB2: data_out = 8'h9;
                    16'h3BB3: data_out = 8'h8;
                    16'h3BB4: data_out = 8'h7;
                    16'h3BB5: data_out = 8'h6;
                    16'h3BB6: data_out = 8'h5;
                    16'h3BB7: data_out = 8'h4;
                    16'h3BB8: data_out = 8'h3;
                    16'h3BB9: data_out = 8'h2;
                    16'h3BBA: data_out = 8'h1;
                    16'h3BBB: data_out = 8'h0;
                    16'h3BBC: data_out = 8'h81;
                    16'h3BBD: data_out = 8'h82;
                    16'h3BBE: data_out = 8'h83;
                    16'h3BBF: data_out = 8'h84;
                    16'h3BC0: data_out = 8'h85;
                    16'h3BC1: data_out = 8'h86;
                    16'h3BC2: data_out = 8'h87;
                    16'h3BC3: data_out = 8'h88;
                    16'h3BC4: data_out = 8'h89;
                    16'h3BC5: data_out = 8'h8A;
                    16'h3BC6: data_out = 8'h8B;
                    16'h3BC7: data_out = 8'h8C;
                    16'h3BC8: data_out = 8'h8D;
                    16'h3BC9: data_out = 8'h8E;
                    16'h3BCA: data_out = 8'h8F;
                    16'h3BCB: data_out = 8'h90;
                    16'h3BCC: data_out = 8'h91;
                    16'h3BCD: data_out = 8'h92;
                    16'h3BCE: data_out = 8'h93;
                    16'h3BCF: data_out = 8'h94;
                    16'h3BD0: data_out = 8'h95;
                    16'h3BD1: data_out = 8'h96;
                    16'h3BD2: data_out = 8'h97;
                    16'h3BD3: data_out = 8'h98;
                    16'h3BD4: data_out = 8'h99;
                    16'h3BD5: data_out = 8'h9A;
                    16'h3BD6: data_out = 8'h9B;
                    16'h3BD7: data_out = 8'h9C;
                    16'h3BD8: data_out = 8'h9D;
                    16'h3BD9: data_out = 8'h9E;
                    16'h3BDA: data_out = 8'h9F;
                    16'h3BDB: data_out = 8'hA0;
                    16'h3BDC: data_out = 8'hA1;
                    16'h3BDD: data_out = 8'hA2;
                    16'h3BDE: data_out = 8'hA3;
                    16'h3BDF: data_out = 8'hA4;
                    16'h3BE0: data_out = 8'hA5;
                    16'h3BE1: data_out = 8'hA6;
                    16'h3BE2: data_out = 8'hA7;
                    16'h3BE3: data_out = 8'hA8;
                    16'h3BE4: data_out = 8'hA9;
                    16'h3BE5: data_out = 8'hAA;
                    16'h3BE6: data_out = 8'hAB;
                    16'h3BE7: data_out = 8'hAC;
                    16'h3BE8: data_out = 8'hAD;
                    16'h3BE9: data_out = 8'hAE;
                    16'h3BEA: data_out = 8'hAF;
                    16'h3BEB: data_out = 8'hB0;
                    16'h3BEC: data_out = 8'hB1;
                    16'h3BED: data_out = 8'hB2;
                    16'h3BEE: data_out = 8'hB3;
                    16'h3BEF: data_out = 8'hB4;
                    16'h3BF0: data_out = 8'hB5;
                    16'h3BF1: data_out = 8'hB6;
                    16'h3BF2: data_out = 8'hB7;
                    16'h3BF3: data_out = 8'hB8;
                    16'h3BF4: data_out = 8'hB9;
                    16'h3BF5: data_out = 8'hBA;
                    16'h3BF6: data_out = 8'hBB;
                    16'h3BF7: data_out = 8'hBC;
                    16'h3BF8: data_out = 8'hBD;
                    16'h3BF9: data_out = 8'hBE;
                    16'h3BFA: data_out = 8'hBF;
                    16'h3BFB: data_out = 8'hC0;
                    16'h3BFC: data_out = 8'hC1;
                    16'h3BFD: data_out = 8'hC2;
                    16'h3BFE: data_out = 8'hC3;
                    16'h3BFF: data_out = 8'hC4;
                    16'h3C00: data_out = 8'h3C;
                    16'h3C01: data_out = 8'h3D;
                    16'h3C02: data_out = 8'h3E;
                    16'h3C03: data_out = 8'h3F;
                    16'h3C04: data_out = 8'h40;
                    16'h3C05: data_out = 8'h41;
                    16'h3C06: data_out = 8'h42;
                    16'h3C07: data_out = 8'h43;
                    16'h3C08: data_out = 8'h44;
                    16'h3C09: data_out = 8'h45;
                    16'h3C0A: data_out = 8'h46;
                    16'h3C0B: data_out = 8'h47;
                    16'h3C0C: data_out = 8'h48;
                    16'h3C0D: data_out = 8'h49;
                    16'h3C0E: data_out = 8'h4A;
                    16'h3C0F: data_out = 8'h4B;
                    16'h3C10: data_out = 8'h4C;
                    16'h3C11: data_out = 8'h4D;
                    16'h3C12: data_out = 8'h4E;
                    16'h3C13: data_out = 8'h4F;
                    16'h3C14: data_out = 8'h50;
                    16'h3C15: data_out = 8'h51;
                    16'h3C16: data_out = 8'h52;
                    16'h3C17: data_out = 8'h53;
                    16'h3C18: data_out = 8'h54;
                    16'h3C19: data_out = 8'h55;
                    16'h3C1A: data_out = 8'h56;
                    16'h3C1B: data_out = 8'h57;
                    16'h3C1C: data_out = 8'h58;
                    16'h3C1D: data_out = 8'h59;
                    16'h3C1E: data_out = 8'h5A;
                    16'h3C1F: data_out = 8'h5B;
                    16'h3C20: data_out = 8'h5C;
                    16'h3C21: data_out = 8'h5D;
                    16'h3C22: data_out = 8'h5E;
                    16'h3C23: data_out = 8'h5F;
                    16'h3C24: data_out = 8'h60;
                    16'h3C25: data_out = 8'h61;
                    16'h3C26: data_out = 8'h62;
                    16'h3C27: data_out = 8'h63;
                    16'h3C28: data_out = 8'h64;
                    16'h3C29: data_out = 8'h65;
                    16'h3C2A: data_out = 8'h66;
                    16'h3C2B: data_out = 8'h67;
                    16'h3C2C: data_out = 8'h68;
                    16'h3C2D: data_out = 8'h69;
                    16'h3C2E: data_out = 8'h6A;
                    16'h3C2F: data_out = 8'h6B;
                    16'h3C30: data_out = 8'h6C;
                    16'h3C31: data_out = 8'h6D;
                    16'h3C32: data_out = 8'h6E;
                    16'h3C33: data_out = 8'h6F;
                    16'h3C34: data_out = 8'h70;
                    16'h3C35: data_out = 8'h71;
                    16'h3C36: data_out = 8'h72;
                    16'h3C37: data_out = 8'h73;
                    16'h3C38: data_out = 8'h74;
                    16'h3C39: data_out = 8'h75;
                    16'h3C3A: data_out = 8'h76;
                    16'h3C3B: data_out = 8'h77;
                    16'h3C3C: data_out = 8'h78;
                    16'h3C3D: data_out = 8'h79;
                    16'h3C3E: data_out = 8'h7A;
                    16'h3C3F: data_out = 8'h7B;
                    16'h3C40: data_out = 8'h7C;
                    16'h3C41: data_out = 8'h7D;
                    16'h3C42: data_out = 8'h7E;
                    16'h3C43: data_out = 8'h7F;
                    16'h3C44: data_out = 8'h80;
                    16'h3C45: data_out = 8'h81;
                    16'h3C46: data_out = 8'h82;
                    16'h3C47: data_out = 8'h83;
                    16'h3C48: data_out = 8'h84;
                    16'h3C49: data_out = 8'h85;
                    16'h3C4A: data_out = 8'h86;
                    16'h3C4B: data_out = 8'h87;
                    16'h3C4C: data_out = 8'h88;
                    16'h3C4D: data_out = 8'h89;
                    16'h3C4E: data_out = 8'h8A;
                    16'h3C4F: data_out = 8'h8B;
                    16'h3C50: data_out = 8'h8C;
                    16'h3C51: data_out = 8'h8D;
                    16'h3C52: data_out = 8'h8E;
                    16'h3C53: data_out = 8'h8F;
                    16'h3C54: data_out = 8'h90;
                    16'h3C55: data_out = 8'h91;
                    16'h3C56: data_out = 8'h92;
                    16'h3C57: data_out = 8'h93;
                    16'h3C58: data_out = 8'h94;
                    16'h3C59: data_out = 8'h95;
                    16'h3C5A: data_out = 8'h96;
                    16'h3C5B: data_out = 8'h97;
                    16'h3C5C: data_out = 8'h98;
                    16'h3C5D: data_out = 8'h99;
                    16'h3C5E: data_out = 8'h9A;
                    16'h3C5F: data_out = 8'h9B;
                    16'h3C60: data_out = 8'h9C;
                    16'h3C61: data_out = 8'h9D;
                    16'h3C62: data_out = 8'h9E;
                    16'h3C63: data_out = 8'h9F;
                    16'h3C64: data_out = 8'hA0;
                    16'h3C65: data_out = 8'hA1;
                    16'h3C66: data_out = 8'hA2;
                    16'h3C67: data_out = 8'hA3;
                    16'h3C68: data_out = 8'hA4;
                    16'h3C69: data_out = 8'hA5;
                    16'h3C6A: data_out = 8'hA6;
                    16'h3C6B: data_out = 8'hA7;
                    16'h3C6C: data_out = 8'hA8;
                    16'h3C6D: data_out = 8'hA9;
                    16'h3C6E: data_out = 8'hAA;
                    16'h3C6F: data_out = 8'hAB;
                    16'h3C70: data_out = 8'hAC;
                    16'h3C71: data_out = 8'hAD;
                    16'h3C72: data_out = 8'hAE;
                    16'h3C73: data_out = 8'hAF;
                    16'h3C74: data_out = 8'hB0;
                    16'h3C75: data_out = 8'hB1;
                    16'h3C76: data_out = 8'hB2;
                    16'h3C77: data_out = 8'hB3;
                    16'h3C78: data_out = 8'hB4;
                    16'h3C79: data_out = 8'hB5;
                    16'h3C7A: data_out = 8'hB6;
                    16'h3C7B: data_out = 8'hB7;
                    16'h3C7C: data_out = 8'hB8;
                    16'h3C7D: data_out = 8'hB9;
                    16'h3C7E: data_out = 8'hBA;
                    16'h3C7F: data_out = 8'hBB;
                    16'h3C80: data_out = 8'h3C;
                    16'h3C81: data_out = 8'h3B;
                    16'h3C82: data_out = 8'h3A;
                    16'h3C83: data_out = 8'h39;
                    16'h3C84: data_out = 8'h38;
                    16'h3C85: data_out = 8'h37;
                    16'h3C86: data_out = 8'h36;
                    16'h3C87: data_out = 8'h35;
                    16'h3C88: data_out = 8'h34;
                    16'h3C89: data_out = 8'h33;
                    16'h3C8A: data_out = 8'h32;
                    16'h3C8B: data_out = 8'h31;
                    16'h3C8C: data_out = 8'h30;
                    16'h3C8D: data_out = 8'h2F;
                    16'h3C8E: data_out = 8'h2E;
                    16'h3C8F: data_out = 8'h2D;
                    16'h3C90: data_out = 8'h2C;
                    16'h3C91: data_out = 8'h2B;
                    16'h3C92: data_out = 8'h2A;
                    16'h3C93: data_out = 8'h29;
                    16'h3C94: data_out = 8'h28;
                    16'h3C95: data_out = 8'h27;
                    16'h3C96: data_out = 8'h26;
                    16'h3C97: data_out = 8'h25;
                    16'h3C98: data_out = 8'h24;
                    16'h3C99: data_out = 8'h23;
                    16'h3C9A: data_out = 8'h22;
                    16'h3C9B: data_out = 8'h21;
                    16'h3C9C: data_out = 8'h20;
                    16'h3C9D: data_out = 8'h1F;
                    16'h3C9E: data_out = 8'h1E;
                    16'h3C9F: data_out = 8'h1D;
                    16'h3CA0: data_out = 8'h1C;
                    16'h3CA1: data_out = 8'h1B;
                    16'h3CA2: data_out = 8'h1A;
                    16'h3CA3: data_out = 8'h19;
                    16'h3CA4: data_out = 8'h18;
                    16'h3CA5: data_out = 8'h17;
                    16'h3CA6: data_out = 8'h16;
                    16'h3CA7: data_out = 8'h15;
                    16'h3CA8: data_out = 8'h14;
                    16'h3CA9: data_out = 8'h13;
                    16'h3CAA: data_out = 8'h12;
                    16'h3CAB: data_out = 8'h11;
                    16'h3CAC: data_out = 8'h10;
                    16'h3CAD: data_out = 8'hF;
                    16'h3CAE: data_out = 8'hE;
                    16'h3CAF: data_out = 8'hD;
                    16'h3CB0: data_out = 8'hC;
                    16'h3CB1: data_out = 8'hB;
                    16'h3CB2: data_out = 8'hA;
                    16'h3CB3: data_out = 8'h9;
                    16'h3CB4: data_out = 8'h8;
                    16'h3CB5: data_out = 8'h7;
                    16'h3CB6: data_out = 8'h6;
                    16'h3CB7: data_out = 8'h5;
                    16'h3CB8: data_out = 8'h4;
                    16'h3CB9: data_out = 8'h3;
                    16'h3CBA: data_out = 8'h2;
                    16'h3CBB: data_out = 8'h1;
                    16'h3CBC: data_out = 8'h0;
                    16'h3CBD: data_out = 8'h81;
                    16'h3CBE: data_out = 8'h82;
                    16'h3CBF: data_out = 8'h83;
                    16'h3CC0: data_out = 8'h84;
                    16'h3CC1: data_out = 8'h85;
                    16'h3CC2: data_out = 8'h86;
                    16'h3CC3: data_out = 8'h87;
                    16'h3CC4: data_out = 8'h88;
                    16'h3CC5: data_out = 8'h89;
                    16'h3CC6: data_out = 8'h8A;
                    16'h3CC7: data_out = 8'h8B;
                    16'h3CC8: data_out = 8'h8C;
                    16'h3CC9: data_out = 8'h8D;
                    16'h3CCA: data_out = 8'h8E;
                    16'h3CCB: data_out = 8'h8F;
                    16'h3CCC: data_out = 8'h90;
                    16'h3CCD: data_out = 8'h91;
                    16'h3CCE: data_out = 8'h92;
                    16'h3CCF: data_out = 8'h93;
                    16'h3CD0: data_out = 8'h94;
                    16'h3CD1: data_out = 8'h95;
                    16'h3CD2: data_out = 8'h96;
                    16'h3CD3: data_out = 8'h97;
                    16'h3CD4: data_out = 8'h98;
                    16'h3CD5: data_out = 8'h99;
                    16'h3CD6: data_out = 8'h9A;
                    16'h3CD7: data_out = 8'h9B;
                    16'h3CD8: data_out = 8'h9C;
                    16'h3CD9: data_out = 8'h9D;
                    16'h3CDA: data_out = 8'h9E;
                    16'h3CDB: data_out = 8'h9F;
                    16'h3CDC: data_out = 8'hA0;
                    16'h3CDD: data_out = 8'hA1;
                    16'h3CDE: data_out = 8'hA2;
                    16'h3CDF: data_out = 8'hA3;
                    16'h3CE0: data_out = 8'hA4;
                    16'h3CE1: data_out = 8'hA5;
                    16'h3CE2: data_out = 8'hA6;
                    16'h3CE3: data_out = 8'hA7;
                    16'h3CE4: data_out = 8'hA8;
                    16'h3CE5: data_out = 8'hA9;
                    16'h3CE6: data_out = 8'hAA;
                    16'h3CE7: data_out = 8'hAB;
                    16'h3CE8: data_out = 8'hAC;
                    16'h3CE9: data_out = 8'hAD;
                    16'h3CEA: data_out = 8'hAE;
                    16'h3CEB: data_out = 8'hAF;
                    16'h3CEC: data_out = 8'hB0;
                    16'h3CED: data_out = 8'hB1;
                    16'h3CEE: data_out = 8'hB2;
                    16'h3CEF: data_out = 8'hB3;
                    16'h3CF0: data_out = 8'hB4;
                    16'h3CF1: data_out = 8'hB5;
                    16'h3CF2: data_out = 8'hB6;
                    16'h3CF3: data_out = 8'hB7;
                    16'h3CF4: data_out = 8'hB8;
                    16'h3CF5: data_out = 8'hB9;
                    16'h3CF6: data_out = 8'hBA;
                    16'h3CF7: data_out = 8'hBB;
                    16'h3CF8: data_out = 8'hBC;
                    16'h3CF9: data_out = 8'hBD;
                    16'h3CFA: data_out = 8'hBE;
                    16'h3CFB: data_out = 8'hBF;
                    16'h3CFC: data_out = 8'hC0;
                    16'h3CFD: data_out = 8'hC1;
                    16'h3CFE: data_out = 8'hC2;
                    16'h3CFF: data_out = 8'hC3;
                    16'h3D00: data_out = 8'h3D;
                    16'h3D01: data_out = 8'h3E;
                    16'h3D02: data_out = 8'h3F;
                    16'h3D03: data_out = 8'h40;
                    16'h3D04: data_out = 8'h41;
                    16'h3D05: data_out = 8'h42;
                    16'h3D06: data_out = 8'h43;
                    16'h3D07: data_out = 8'h44;
                    16'h3D08: data_out = 8'h45;
                    16'h3D09: data_out = 8'h46;
                    16'h3D0A: data_out = 8'h47;
                    16'h3D0B: data_out = 8'h48;
                    16'h3D0C: data_out = 8'h49;
                    16'h3D0D: data_out = 8'h4A;
                    16'h3D0E: data_out = 8'h4B;
                    16'h3D0F: data_out = 8'h4C;
                    16'h3D10: data_out = 8'h4D;
                    16'h3D11: data_out = 8'h4E;
                    16'h3D12: data_out = 8'h4F;
                    16'h3D13: data_out = 8'h50;
                    16'h3D14: data_out = 8'h51;
                    16'h3D15: data_out = 8'h52;
                    16'h3D16: data_out = 8'h53;
                    16'h3D17: data_out = 8'h54;
                    16'h3D18: data_out = 8'h55;
                    16'h3D19: data_out = 8'h56;
                    16'h3D1A: data_out = 8'h57;
                    16'h3D1B: data_out = 8'h58;
                    16'h3D1C: data_out = 8'h59;
                    16'h3D1D: data_out = 8'h5A;
                    16'h3D1E: data_out = 8'h5B;
                    16'h3D1F: data_out = 8'h5C;
                    16'h3D20: data_out = 8'h5D;
                    16'h3D21: data_out = 8'h5E;
                    16'h3D22: data_out = 8'h5F;
                    16'h3D23: data_out = 8'h60;
                    16'h3D24: data_out = 8'h61;
                    16'h3D25: data_out = 8'h62;
                    16'h3D26: data_out = 8'h63;
                    16'h3D27: data_out = 8'h64;
                    16'h3D28: data_out = 8'h65;
                    16'h3D29: data_out = 8'h66;
                    16'h3D2A: data_out = 8'h67;
                    16'h3D2B: data_out = 8'h68;
                    16'h3D2C: data_out = 8'h69;
                    16'h3D2D: data_out = 8'h6A;
                    16'h3D2E: data_out = 8'h6B;
                    16'h3D2F: data_out = 8'h6C;
                    16'h3D30: data_out = 8'h6D;
                    16'h3D31: data_out = 8'h6E;
                    16'h3D32: data_out = 8'h6F;
                    16'h3D33: data_out = 8'h70;
                    16'h3D34: data_out = 8'h71;
                    16'h3D35: data_out = 8'h72;
                    16'h3D36: data_out = 8'h73;
                    16'h3D37: data_out = 8'h74;
                    16'h3D38: data_out = 8'h75;
                    16'h3D39: data_out = 8'h76;
                    16'h3D3A: data_out = 8'h77;
                    16'h3D3B: data_out = 8'h78;
                    16'h3D3C: data_out = 8'h79;
                    16'h3D3D: data_out = 8'h7A;
                    16'h3D3E: data_out = 8'h7B;
                    16'h3D3F: data_out = 8'h7C;
                    16'h3D40: data_out = 8'h7D;
                    16'h3D41: data_out = 8'h7E;
                    16'h3D42: data_out = 8'h7F;
                    16'h3D43: data_out = 8'h80;
                    16'h3D44: data_out = 8'h81;
                    16'h3D45: data_out = 8'h82;
                    16'h3D46: data_out = 8'h83;
                    16'h3D47: data_out = 8'h84;
                    16'h3D48: data_out = 8'h85;
                    16'h3D49: data_out = 8'h86;
                    16'h3D4A: data_out = 8'h87;
                    16'h3D4B: data_out = 8'h88;
                    16'h3D4C: data_out = 8'h89;
                    16'h3D4D: data_out = 8'h8A;
                    16'h3D4E: data_out = 8'h8B;
                    16'h3D4F: data_out = 8'h8C;
                    16'h3D50: data_out = 8'h8D;
                    16'h3D51: data_out = 8'h8E;
                    16'h3D52: data_out = 8'h8F;
                    16'h3D53: data_out = 8'h90;
                    16'h3D54: data_out = 8'h91;
                    16'h3D55: data_out = 8'h92;
                    16'h3D56: data_out = 8'h93;
                    16'h3D57: data_out = 8'h94;
                    16'h3D58: data_out = 8'h95;
                    16'h3D59: data_out = 8'h96;
                    16'h3D5A: data_out = 8'h97;
                    16'h3D5B: data_out = 8'h98;
                    16'h3D5C: data_out = 8'h99;
                    16'h3D5D: data_out = 8'h9A;
                    16'h3D5E: data_out = 8'h9B;
                    16'h3D5F: data_out = 8'h9C;
                    16'h3D60: data_out = 8'h9D;
                    16'h3D61: data_out = 8'h9E;
                    16'h3D62: data_out = 8'h9F;
                    16'h3D63: data_out = 8'hA0;
                    16'h3D64: data_out = 8'hA1;
                    16'h3D65: data_out = 8'hA2;
                    16'h3D66: data_out = 8'hA3;
                    16'h3D67: data_out = 8'hA4;
                    16'h3D68: data_out = 8'hA5;
                    16'h3D69: data_out = 8'hA6;
                    16'h3D6A: data_out = 8'hA7;
                    16'h3D6B: data_out = 8'hA8;
                    16'h3D6C: data_out = 8'hA9;
                    16'h3D6D: data_out = 8'hAA;
                    16'h3D6E: data_out = 8'hAB;
                    16'h3D6F: data_out = 8'hAC;
                    16'h3D70: data_out = 8'hAD;
                    16'h3D71: data_out = 8'hAE;
                    16'h3D72: data_out = 8'hAF;
                    16'h3D73: data_out = 8'hB0;
                    16'h3D74: data_out = 8'hB1;
                    16'h3D75: data_out = 8'hB2;
                    16'h3D76: data_out = 8'hB3;
                    16'h3D77: data_out = 8'hB4;
                    16'h3D78: data_out = 8'hB5;
                    16'h3D79: data_out = 8'hB6;
                    16'h3D7A: data_out = 8'hB7;
                    16'h3D7B: data_out = 8'hB8;
                    16'h3D7C: data_out = 8'hB9;
                    16'h3D7D: data_out = 8'hBA;
                    16'h3D7E: data_out = 8'hBB;
                    16'h3D7F: data_out = 8'hBC;
                    16'h3D80: data_out = 8'h3D;
                    16'h3D81: data_out = 8'h3C;
                    16'h3D82: data_out = 8'h3B;
                    16'h3D83: data_out = 8'h3A;
                    16'h3D84: data_out = 8'h39;
                    16'h3D85: data_out = 8'h38;
                    16'h3D86: data_out = 8'h37;
                    16'h3D87: data_out = 8'h36;
                    16'h3D88: data_out = 8'h35;
                    16'h3D89: data_out = 8'h34;
                    16'h3D8A: data_out = 8'h33;
                    16'h3D8B: data_out = 8'h32;
                    16'h3D8C: data_out = 8'h31;
                    16'h3D8D: data_out = 8'h30;
                    16'h3D8E: data_out = 8'h2F;
                    16'h3D8F: data_out = 8'h2E;
                    16'h3D90: data_out = 8'h2D;
                    16'h3D91: data_out = 8'h2C;
                    16'h3D92: data_out = 8'h2B;
                    16'h3D93: data_out = 8'h2A;
                    16'h3D94: data_out = 8'h29;
                    16'h3D95: data_out = 8'h28;
                    16'h3D96: data_out = 8'h27;
                    16'h3D97: data_out = 8'h26;
                    16'h3D98: data_out = 8'h25;
                    16'h3D99: data_out = 8'h24;
                    16'h3D9A: data_out = 8'h23;
                    16'h3D9B: data_out = 8'h22;
                    16'h3D9C: data_out = 8'h21;
                    16'h3D9D: data_out = 8'h20;
                    16'h3D9E: data_out = 8'h1F;
                    16'h3D9F: data_out = 8'h1E;
                    16'h3DA0: data_out = 8'h1D;
                    16'h3DA1: data_out = 8'h1C;
                    16'h3DA2: data_out = 8'h1B;
                    16'h3DA3: data_out = 8'h1A;
                    16'h3DA4: data_out = 8'h19;
                    16'h3DA5: data_out = 8'h18;
                    16'h3DA6: data_out = 8'h17;
                    16'h3DA7: data_out = 8'h16;
                    16'h3DA8: data_out = 8'h15;
                    16'h3DA9: data_out = 8'h14;
                    16'h3DAA: data_out = 8'h13;
                    16'h3DAB: data_out = 8'h12;
                    16'h3DAC: data_out = 8'h11;
                    16'h3DAD: data_out = 8'h10;
                    16'h3DAE: data_out = 8'hF;
                    16'h3DAF: data_out = 8'hE;
                    16'h3DB0: data_out = 8'hD;
                    16'h3DB1: data_out = 8'hC;
                    16'h3DB2: data_out = 8'hB;
                    16'h3DB3: data_out = 8'hA;
                    16'h3DB4: data_out = 8'h9;
                    16'h3DB5: data_out = 8'h8;
                    16'h3DB6: data_out = 8'h7;
                    16'h3DB7: data_out = 8'h6;
                    16'h3DB8: data_out = 8'h5;
                    16'h3DB9: data_out = 8'h4;
                    16'h3DBA: data_out = 8'h3;
                    16'h3DBB: data_out = 8'h2;
                    16'h3DBC: data_out = 8'h1;
                    16'h3DBD: data_out = 8'h0;
                    16'h3DBE: data_out = 8'h81;
                    16'h3DBF: data_out = 8'h82;
                    16'h3DC0: data_out = 8'h83;
                    16'h3DC1: data_out = 8'h84;
                    16'h3DC2: data_out = 8'h85;
                    16'h3DC3: data_out = 8'h86;
                    16'h3DC4: data_out = 8'h87;
                    16'h3DC5: data_out = 8'h88;
                    16'h3DC6: data_out = 8'h89;
                    16'h3DC7: data_out = 8'h8A;
                    16'h3DC8: data_out = 8'h8B;
                    16'h3DC9: data_out = 8'h8C;
                    16'h3DCA: data_out = 8'h8D;
                    16'h3DCB: data_out = 8'h8E;
                    16'h3DCC: data_out = 8'h8F;
                    16'h3DCD: data_out = 8'h90;
                    16'h3DCE: data_out = 8'h91;
                    16'h3DCF: data_out = 8'h92;
                    16'h3DD0: data_out = 8'h93;
                    16'h3DD1: data_out = 8'h94;
                    16'h3DD2: data_out = 8'h95;
                    16'h3DD3: data_out = 8'h96;
                    16'h3DD4: data_out = 8'h97;
                    16'h3DD5: data_out = 8'h98;
                    16'h3DD6: data_out = 8'h99;
                    16'h3DD7: data_out = 8'h9A;
                    16'h3DD8: data_out = 8'h9B;
                    16'h3DD9: data_out = 8'h9C;
                    16'h3DDA: data_out = 8'h9D;
                    16'h3DDB: data_out = 8'h9E;
                    16'h3DDC: data_out = 8'h9F;
                    16'h3DDD: data_out = 8'hA0;
                    16'h3DDE: data_out = 8'hA1;
                    16'h3DDF: data_out = 8'hA2;
                    16'h3DE0: data_out = 8'hA3;
                    16'h3DE1: data_out = 8'hA4;
                    16'h3DE2: data_out = 8'hA5;
                    16'h3DE3: data_out = 8'hA6;
                    16'h3DE4: data_out = 8'hA7;
                    16'h3DE5: data_out = 8'hA8;
                    16'h3DE6: data_out = 8'hA9;
                    16'h3DE7: data_out = 8'hAA;
                    16'h3DE8: data_out = 8'hAB;
                    16'h3DE9: data_out = 8'hAC;
                    16'h3DEA: data_out = 8'hAD;
                    16'h3DEB: data_out = 8'hAE;
                    16'h3DEC: data_out = 8'hAF;
                    16'h3DED: data_out = 8'hB0;
                    16'h3DEE: data_out = 8'hB1;
                    16'h3DEF: data_out = 8'hB2;
                    16'h3DF0: data_out = 8'hB3;
                    16'h3DF1: data_out = 8'hB4;
                    16'h3DF2: data_out = 8'hB5;
                    16'h3DF3: data_out = 8'hB6;
                    16'h3DF4: data_out = 8'hB7;
                    16'h3DF5: data_out = 8'hB8;
                    16'h3DF6: data_out = 8'hB9;
                    16'h3DF7: data_out = 8'hBA;
                    16'h3DF8: data_out = 8'hBB;
                    16'h3DF9: data_out = 8'hBC;
                    16'h3DFA: data_out = 8'hBD;
                    16'h3DFB: data_out = 8'hBE;
                    16'h3DFC: data_out = 8'hBF;
                    16'h3DFD: data_out = 8'hC0;
                    16'h3DFE: data_out = 8'hC1;
                    16'h3DFF: data_out = 8'hC2;
                    16'h3E00: data_out = 8'h3E;
                    16'h3E01: data_out = 8'h3F;
                    16'h3E02: data_out = 8'h40;
                    16'h3E03: data_out = 8'h41;
                    16'h3E04: data_out = 8'h42;
                    16'h3E05: data_out = 8'h43;
                    16'h3E06: data_out = 8'h44;
                    16'h3E07: data_out = 8'h45;
                    16'h3E08: data_out = 8'h46;
                    16'h3E09: data_out = 8'h47;
                    16'h3E0A: data_out = 8'h48;
                    16'h3E0B: data_out = 8'h49;
                    16'h3E0C: data_out = 8'h4A;
                    16'h3E0D: data_out = 8'h4B;
                    16'h3E0E: data_out = 8'h4C;
                    16'h3E0F: data_out = 8'h4D;
                    16'h3E10: data_out = 8'h4E;
                    16'h3E11: data_out = 8'h4F;
                    16'h3E12: data_out = 8'h50;
                    16'h3E13: data_out = 8'h51;
                    16'h3E14: data_out = 8'h52;
                    16'h3E15: data_out = 8'h53;
                    16'h3E16: data_out = 8'h54;
                    16'h3E17: data_out = 8'h55;
                    16'h3E18: data_out = 8'h56;
                    16'h3E19: data_out = 8'h57;
                    16'h3E1A: data_out = 8'h58;
                    16'h3E1B: data_out = 8'h59;
                    16'h3E1C: data_out = 8'h5A;
                    16'h3E1D: data_out = 8'h5B;
                    16'h3E1E: data_out = 8'h5C;
                    16'h3E1F: data_out = 8'h5D;
                    16'h3E20: data_out = 8'h5E;
                    16'h3E21: data_out = 8'h5F;
                    16'h3E22: data_out = 8'h60;
                    16'h3E23: data_out = 8'h61;
                    16'h3E24: data_out = 8'h62;
                    16'h3E25: data_out = 8'h63;
                    16'h3E26: data_out = 8'h64;
                    16'h3E27: data_out = 8'h65;
                    16'h3E28: data_out = 8'h66;
                    16'h3E29: data_out = 8'h67;
                    16'h3E2A: data_out = 8'h68;
                    16'h3E2B: data_out = 8'h69;
                    16'h3E2C: data_out = 8'h6A;
                    16'h3E2D: data_out = 8'h6B;
                    16'h3E2E: data_out = 8'h6C;
                    16'h3E2F: data_out = 8'h6D;
                    16'h3E30: data_out = 8'h6E;
                    16'h3E31: data_out = 8'h6F;
                    16'h3E32: data_out = 8'h70;
                    16'h3E33: data_out = 8'h71;
                    16'h3E34: data_out = 8'h72;
                    16'h3E35: data_out = 8'h73;
                    16'h3E36: data_out = 8'h74;
                    16'h3E37: data_out = 8'h75;
                    16'h3E38: data_out = 8'h76;
                    16'h3E39: data_out = 8'h77;
                    16'h3E3A: data_out = 8'h78;
                    16'h3E3B: data_out = 8'h79;
                    16'h3E3C: data_out = 8'h7A;
                    16'h3E3D: data_out = 8'h7B;
                    16'h3E3E: data_out = 8'h7C;
                    16'h3E3F: data_out = 8'h7D;
                    16'h3E40: data_out = 8'h7E;
                    16'h3E41: data_out = 8'h7F;
                    16'h3E42: data_out = 8'h80;
                    16'h3E43: data_out = 8'h81;
                    16'h3E44: data_out = 8'h82;
                    16'h3E45: data_out = 8'h83;
                    16'h3E46: data_out = 8'h84;
                    16'h3E47: data_out = 8'h85;
                    16'h3E48: data_out = 8'h86;
                    16'h3E49: data_out = 8'h87;
                    16'h3E4A: data_out = 8'h88;
                    16'h3E4B: data_out = 8'h89;
                    16'h3E4C: data_out = 8'h8A;
                    16'h3E4D: data_out = 8'h8B;
                    16'h3E4E: data_out = 8'h8C;
                    16'h3E4F: data_out = 8'h8D;
                    16'h3E50: data_out = 8'h8E;
                    16'h3E51: data_out = 8'h8F;
                    16'h3E52: data_out = 8'h90;
                    16'h3E53: data_out = 8'h91;
                    16'h3E54: data_out = 8'h92;
                    16'h3E55: data_out = 8'h93;
                    16'h3E56: data_out = 8'h94;
                    16'h3E57: data_out = 8'h95;
                    16'h3E58: data_out = 8'h96;
                    16'h3E59: data_out = 8'h97;
                    16'h3E5A: data_out = 8'h98;
                    16'h3E5B: data_out = 8'h99;
                    16'h3E5C: data_out = 8'h9A;
                    16'h3E5D: data_out = 8'h9B;
                    16'h3E5E: data_out = 8'h9C;
                    16'h3E5F: data_out = 8'h9D;
                    16'h3E60: data_out = 8'h9E;
                    16'h3E61: data_out = 8'h9F;
                    16'h3E62: data_out = 8'hA0;
                    16'h3E63: data_out = 8'hA1;
                    16'h3E64: data_out = 8'hA2;
                    16'h3E65: data_out = 8'hA3;
                    16'h3E66: data_out = 8'hA4;
                    16'h3E67: data_out = 8'hA5;
                    16'h3E68: data_out = 8'hA6;
                    16'h3E69: data_out = 8'hA7;
                    16'h3E6A: data_out = 8'hA8;
                    16'h3E6B: data_out = 8'hA9;
                    16'h3E6C: data_out = 8'hAA;
                    16'h3E6D: data_out = 8'hAB;
                    16'h3E6E: data_out = 8'hAC;
                    16'h3E6F: data_out = 8'hAD;
                    16'h3E70: data_out = 8'hAE;
                    16'h3E71: data_out = 8'hAF;
                    16'h3E72: data_out = 8'hB0;
                    16'h3E73: data_out = 8'hB1;
                    16'h3E74: data_out = 8'hB2;
                    16'h3E75: data_out = 8'hB3;
                    16'h3E76: data_out = 8'hB4;
                    16'h3E77: data_out = 8'hB5;
                    16'h3E78: data_out = 8'hB6;
                    16'h3E79: data_out = 8'hB7;
                    16'h3E7A: data_out = 8'hB8;
                    16'h3E7B: data_out = 8'hB9;
                    16'h3E7C: data_out = 8'hBA;
                    16'h3E7D: data_out = 8'hBB;
                    16'h3E7E: data_out = 8'hBC;
                    16'h3E7F: data_out = 8'hBD;
                    16'h3E80: data_out = 8'h3E;
                    16'h3E81: data_out = 8'h3D;
                    16'h3E82: data_out = 8'h3C;
                    16'h3E83: data_out = 8'h3B;
                    16'h3E84: data_out = 8'h3A;
                    16'h3E85: data_out = 8'h39;
                    16'h3E86: data_out = 8'h38;
                    16'h3E87: data_out = 8'h37;
                    16'h3E88: data_out = 8'h36;
                    16'h3E89: data_out = 8'h35;
                    16'h3E8A: data_out = 8'h34;
                    16'h3E8B: data_out = 8'h33;
                    16'h3E8C: data_out = 8'h32;
                    16'h3E8D: data_out = 8'h31;
                    16'h3E8E: data_out = 8'h30;
                    16'h3E8F: data_out = 8'h2F;
                    16'h3E90: data_out = 8'h2E;
                    16'h3E91: data_out = 8'h2D;
                    16'h3E92: data_out = 8'h2C;
                    16'h3E93: data_out = 8'h2B;
                    16'h3E94: data_out = 8'h2A;
                    16'h3E95: data_out = 8'h29;
                    16'h3E96: data_out = 8'h28;
                    16'h3E97: data_out = 8'h27;
                    16'h3E98: data_out = 8'h26;
                    16'h3E99: data_out = 8'h25;
                    16'h3E9A: data_out = 8'h24;
                    16'h3E9B: data_out = 8'h23;
                    16'h3E9C: data_out = 8'h22;
                    16'h3E9D: data_out = 8'h21;
                    16'h3E9E: data_out = 8'h20;
                    16'h3E9F: data_out = 8'h1F;
                    16'h3EA0: data_out = 8'h1E;
                    16'h3EA1: data_out = 8'h1D;
                    16'h3EA2: data_out = 8'h1C;
                    16'h3EA3: data_out = 8'h1B;
                    16'h3EA4: data_out = 8'h1A;
                    16'h3EA5: data_out = 8'h19;
                    16'h3EA6: data_out = 8'h18;
                    16'h3EA7: data_out = 8'h17;
                    16'h3EA8: data_out = 8'h16;
                    16'h3EA9: data_out = 8'h15;
                    16'h3EAA: data_out = 8'h14;
                    16'h3EAB: data_out = 8'h13;
                    16'h3EAC: data_out = 8'h12;
                    16'h3EAD: data_out = 8'h11;
                    16'h3EAE: data_out = 8'h10;
                    16'h3EAF: data_out = 8'hF;
                    16'h3EB0: data_out = 8'hE;
                    16'h3EB1: data_out = 8'hD;
                    16'h3EB2: data_out = 8'hC;
                    16'h3EB3: data_out = 8'hB;
                    16'h3EB4: data_out = 8'hA;
                    16'h3EB5: data_out = 8'h9;
                    16'h3EB6: data_out = 8'h8;
                    16'h3EB7: data_out = 8'h7;
                    16'h3EB8: data_out = 8'h6;
                    16'h3EB9: data_out = 8'h5;
                    16'h3EBA: data_out = 8'h4;
                    16'h3EBB: data_out = 8'h3;
                    16'h3EBC: data_out = 8'h2;
                    16'h3EBD: data_out = 8'h1;
                    16'h3EBE: data_out = 8'h0;
                    16'h3EBF: data_out = 8'h81;
                    16'h3EC0: data_out = 8'h82;
                    16'h3EC1: data_out = 8'h83;
                    16'h3EC2: data_out = 8'h84;
                    16'h3EC3: data_out = 8'h85;
                    16'h3EC4: data_out = 8'h86;
                    16'h3EC5: data_out = 8'h87;
                    16'h3EC6: data_out = 8'h88;
                    16'h3EC7: data_out = 8'h89;
                    16'h3EC8: data_out = 8'h8A;
                    16'h3EC9: data_out = 8'h8B;
                    16'h3ECA: data_out = 8'h8C;
                    16'h3ECB: data_out = 8'h8D;
                    16'h3ECC: data_out = 8'h8E;
                    16'h3ECD: data_out = 8'h8F;
                    16'h3ECE: data_out = 8'h90;
                    16'h3ECF: data_out = 8'h91;
                    16'h3ED0: data_out = 8'h92;
                    16'h3ED1: data_out = 8'h93;
                    16'h3ED2: data_out = 8'h94;
                    16'h3ED3: data_out = 8'h95;
                    16'h3ED4: data_out = 8'h96;
                    16'h3ED5: data_out = 8'h97;
                    16'h3ED6: data_out = 8'h98;
                    16'h3ED7: data_out = 8'h99;
                    16'h3ED8: data_out = 8'h9A;
                    16'h3ED9: data_out = 8'h9B;
                    16'h3EDA: data_out = 8'h9C;
                    16'h3EDB: data_out = 8'h9D;
                    16'h3EDC: data_out = 8'h9E;
                    16'h3EDD: data_out = 8'h9F;
                    16'h3EDE: data_out = 8'hA0;
                    16'h3EDF: data_out = 8'hA1;
                    16'h3EE0: data_out = 8'hA2;
                    16'h3EE1: data_out = 8'hA3;
                    16'h3EE2: data_out = 8'hA4;
                    16'h3EE3: data_out = 8'hA5;
                    16'h3EE4: data_out = 8'hA6;
                    16'h3EE5: data_out = 8'hA7;
                    16'h3EE6: data_out = 8'hA8;
                    16'h3EE7: data_out = 8'hA9;
                    16'h3EE8: data_out = 8'hAA;
                    16'h3EE9: data_out = 8'hAB;
                    16'h3EEA: data_out = 8'hAC;
                    16'h3EEB: data_out = 8'hAD;
                    16'h3EEC: data_out = 8'hAE;
                    16'h3EED: data_out = 8'hAF;
                    16'h3EEE: data_out = 8'hB0;
                    16'h3EEF: data_out = 8'hB1;
                    16'h3EF0: data_out = 8'hB2;
                    16'h3EF1: data_out = 8'hB3;
                    16'h3EF2: data_out = 8'hB4;
                    16'h3EF3: data_out = 8'hB5;
                    16'h3EF4: data_out = 8'hB6;
                    16'h3EF5: data_out = 8'hB7;
                    16'h3EF6: data_out = 8'hB8;
                    16'h3EF7: data_out = 8'hB9;
                    16'h3EF8: data_out = 8'hBA;
                    16'h3EF9: data_out = 8'hBB;
                    16'h3EFA: data_out = 8'hBC;
                    16'h3EFB: data_out = 8'hBD;
                    16'h3EFC: data_out = 8'hBE;
                    16'h3EFD: data_out = 8'hBF;
                    16'h3EFE: data_out = 8'hC0;
                    16'h3EFF: data_out = 8'hC1;
                    16'h3F00: data_out = 8'h3F;
                    16'h3F01: data_out = 8'h40;
                    16'h3F02: data_out = 8'h41;
                    16'h3F03: data_out = 8'h42;
                    16'h3F04: data_out = 8'h43;
                    16'h3F05: data_out = 8'h44;
                    16'h3F06: data_out = 8'h45;
                    16'h3F07: data_out = 8'h46;
                    16'h3F08: data_out = 8'h47;
                    16'h3F09: data_out = 8'h48;
                    16'h3F0A: data_out = 8'h49;
                    16'h3F0B: data_out = 8'h4A;
                    16'h3F0C: data_out = 8'h4B;
                    16'h3F0D: data_out = 8'h4C;
                    16'h3F0E: data_out = 8'h4D;
                    16'h3F0F: data_out = 8'h4E;
                    16'h3F10: data_out = 8'h4F;
                    16'h3F11: data_out = 8'h50;
                    16'h3F12: data_out = 8'h51;
                    16'h3F13: data_out = 8'h52;
                    16'h3F14: data_out = 8'h53;
                    16'h3F15: data_out = 8'h54;
                    16'h3F16: data_out = 8'h55;
                    16'h3F17: data_out = 8'h56;
                    16'h3F18: data_out = 8'h57;
                    16'h3F19: data_out = 8'h58;
                    16'h3F1A: data_out = 8'h59;
                    16'h3F1B: data_out = 8'h5A;
                    16'h3F1C: data_out = 8'h5B;
                    16'h3F1D: data_out = 8'h5C;
                    16'h3F1E: data_out = 8'h5D;
                    16'h3F1F: data_out = 8'h5E;
                    16'h3F20: data_out = 8'h5F;
                    16'h3F21: data_out = 8'h60;
                    16'h3F22: data_out = 8'h61;
                    16'h3F23: data_out = 8'h62;
                    16'h3F24: data_out = 8'h63;
                    16'h3F25: data_out = 8'h64;
                    16'h3F26: data_out = 8'h65;
                    16'h3F27: data_out = 8'h66;
                    16'h3F28: data_out = 8'h67;
                    16'h3F29: data_out = 8'h68;
                    16'h3F2A: data_out = 8'h69;
                    16'h3F2B: data_out = 8'h6A;
                    16'h3F2C: data_out = 8'h6B;
                    16'h3F2D: data_out = 8'h6C;
                    16'h3F2E: data_out = 8'h6D;
                    16'h3F2F: data_out = 8'h6E;
                    16'h3F30: data_out = 8'h6F;
                    16'h3F31: data_out = 8'h70;
                    16'h3F32: data_out = 8'h71;
                    16'h3F33: data_out = 8'h72;
                    16'h3F34: data_out = 8'h73;
                    16'h3F35: data_out = 8'h74;
                    16'h3F36: data_out = 8'h75;
                    16'h3F37: data_out = 8'h76;
                    16'h3F38: data_out = 8'h77;
                    16'h3F39: data_out = 8'h78;
                    16'h3F3A: data_out = 8'h79;
                    16'h3F3B: data_out = 8'h7A;
                    16'h3F3C: data_out = 8'h7B;
                    16'h3F3D: data_out = 8'h7C;
                    16'h3F3E: data_out = 8'h7D;
                    16'h3F3F: data_out = 8'h7E;
                    16'h3F40: data_out = 8'h7F;
                    16'h3F41: data_out = 8'h80;
                    16'h3F42: data_out = 8'h81;
                    16'h3F43: data_out = 8'h82;
                    16'h3F44: data_out = 8'h83;
                    16'h3F45: data_out = 8'h84;
                    16'h3F46: data_out = 8'h85;
                    16'h3F47: data_out = 8'h86;
                    16'h3F48: data_out = 8'h87;
                    16'h3F49: data_out = 8'h88;
                    16'h3F4A: data_out = 8'h89;
                    16'h3F4B: data_out = 8'h8A;
                    16'h3F4C: data_out = 8'h8B;
                    16'h3F4D: data_out = 8'h8C;
                    16'h3F4E: data_out = 8'h8D;
                    16'h3F4F: data_out = 8'h8E;
                    16'h3F50: data_out = 8'h8F;
                    16'h3F51: data_out = 8'h90;
                    16'h3F52: data_out = 8'h91;
                    16'h3F53: data_out = 8'h92;
                    16'h3F54: data_out = 8'h93;
                    16'h3F55: data_out = 8'h94;
                    16'h3F56: data_out = 8'h95;
                    16'h3F57: data_out = 8'h96;
                    16'h3F58: data_out = 8'h97;
                    16'h3F59: data_out = 8'h98;
                    16'h3F5A: data_out = 8'h99;
                    16'h3F5B: data_out = 8'h9A;
                    16'h3F5C: data_out = 8'h9B;
                    16'h3F5D: data_out = 8'h9C;
                    16'h3F5E: data_out = 8'h9D;
                    16'h3F5F: data_out = 8'h9E;
                    16'h3F60: data_out = 8'h9F;
                    16'h3F61: data_out = 8'hA0;
                    16'h3F62: data_out = 8'hA1;
                    16'h3F63: data_out = 8'hA2;
                    16'h3F64: data_out = 8'hA3;
                    16'h3F65: data_out = 8'hA4;
                    16'h3F66: data_out = 8'hA5;
                    16'h3F67: data_out = 8'hA6;
                    16'h3F68: data_out = 8'hA7;
                    16'h3F69: data_out = 8'hA8;
                    16'h3F6A: data_out = 8'hA9;
                    16'h3F6B: data_out = 8'hAA;
                    16'h3F6C: data_out = 8'hAB;
                    16'h3F6D: data_out = 8'hAC;
                    16'h3F6E: data_out = 8'hAD;
                    16'h3F6F: data_out = 8'hAE;
                    16'h3F70: data_out = 8'hAF;
                    16'h3F71: data_out = 8'hB0;
                    16'h3F72: data_out = 8'hB1;
                    16'h3F73: data_out = 8'hB2;
                    16'h3F74: data_out = 8'hB3;
                    16'h3F75: data_out = 8'hB4;
                    16'h3F76: data_out = 8'hB5;
                    16'h3F77: data_out = 8'hB6;
                    16'h3F78: data_out = 8'hB7;
                    16'h3F79: data_out = 8'hB8;
                    16'h3F7A: data_out = 8'hB9;
                    16'h3F7B: data_out = 8'hBA;
                    16'h3F7C: data_out = 8'hBB;
                    16'h3F7D: data_out = 8'hBC;
                    16'h3F7E: data_out = 8'hBD;
                    16'h3F7F: data_out = 8'hBE;
                    16'h3F80: data_out = 8'h3F;
                    16'h3F81: data_out = 8'h3E;
                    16'h3F82: data_out = 8'h3D;
                    16'h3F83: data_out = 8'h3C;
                    16'h3F84: data_out = 8'h3B;
                    16'h3F85: data_out = 8'h3A;
                    16'h3F86: data_out = 8'h39;
                    16'h3F87: data_out = 8'h38;
                    16'h3F88: data_out = 8'h37;
                    16'h3F89: data_out = 8'h36;
                    16'h3F8A: data_out = 8'h35;
                    16'h3F8B: data_out = 8'h34;
                    16'h3F8C: data_out = 8'h33;
                    16'h3F8D: data_out = 8'h32;
                    16'h3F8E: data_out = 8'h31;
                    16'h3F8F: data_out = 8'h30;
                    16'h3F90: data_out = 8'h2F;
                    16'h3F91: data_out = 8'h2E;
                    16'h3F92: data_out = 8'h2D;
                    16'h3F93: data_out = 8'h2C;
                    16'h3F94: data_out = 8'h2B;
                    16'h3F95: data_out = 8'h2A;
                    16'h3F96: data_out = 8'h29;
                    16'h3F97: data_out = 8'h28;
                    16'h3F98: data_out = 8'h27;
                    16'h3F99: data_out = 8'h26;
                    16'h3F9A: data_out = 8'h25;
                    16'h3F9B: data_out = 8'h24;
                    16'h3F9C: data_out = 8'h23;
                    16'h3F9D: data_out = 8'h22;
                    16'h3F9E: data_out = 8'h21;
                    16'h3F9F: data_out = 8'h20;
                    16'h3FA0: data_out = 8'h1F;
                    16'h3FA1: data_out = 8'h1E;
                    16'h3FA2: data_out = 8'h1D;
                    16'h3FA3: data_out = 8'h1C;
                    16'h3FA4: data_out = 8'h1B;
                    16'h3FA5: data_out = 8'h1A;
                    16'h3FA6: data_out = 8'h19;
                    16'h3FA7: data_out = 8'h18;
                    16'h3FA8: data_out = 8'h17;
                    16'h3FA9: data_out = 8'h16;
                    16'h3FAA: data_out = 8'h15;
                    16'h3FAB: data_out = 8'h14;
                    16'h3FAC: data_out = 8'h13;
                    16'h3FAD: data_out = 8'h12;
                    16'h3FAE: data_out = 8'h11;
                    16'h3FAF: data_out = 8'h10;
                    16'h3FB0: data_out = 8'hF;
                    16'h3FB1: data_out = 8'hE;
                    16'h3FB2: data_out = 8'hD;
                    16'h3FB3: data_out = 8'hC;
                    16'h3FB4: data_out = 8'hB;
                    16'h3FB5: data_out = 8'hA;
                    16'h3FB6: data_out = 8'h9;
                    16'h3FB7: data_out = 8'h8;
                    16'h3FB8: data_out = 8'h7;
                    16'h3FB9: data_out = 8'h6;
                    16'h3FBA: data_out = 8'h5;
                    16'h3FBB: data_out = 8'h4;
                    16'h3FBC: data_out = 8'h3;
                    16'h3FBD: data_out = 8'h2;
                    16'h3FBE: data_out = 8'h1;
                    16'h3FBF: data_out = 8'h0;
                    16'h3FC0: data_out = 8'h81;
                    16'h3FC1: data_out = 8'h82;
                    16'h3FC2: data_out = 8'h83;
                    16'h3FC3: data_out = 8'h84;
                    16'h3FC4: data_out = 8'h85;
                    16'h3FC5: data_out = 8'h86;
                    16'h3FC6: data_out = 8'h87;
                    16'h3FC7: data_out = 8'h88;
                    16'h3FC8: data_out = 8'h89;
                    16'h3FC9: data_out = 8'h8A;
                    16'h3FCA: data_out = 8'h8B;
                    16'h3FCB: data_out = 8'h8C;
                    16'h3FCC: data_out = 8'h8D;
                    16'h3FCD: data_out = 8'h8E;
                    16'h3FCE: data_out = 8'h8F;
                    16'h3FCF: data_out = 8'h90;
                    16'h3FD0: data_out = 8'h91;
                    16'h3FD1: data_out = 8'h92;
                    16'h3FD2: data_out = 8'h93;
                    16'h3FD3: data_out = 8'h94;
                    16'h3FD4: data_out = 8'h95;
                    16'h3FD5: data_out = 8'h96;
                    16'h3FD6: data_out = 8'h97;
                    16'h3FD7: data_out = 8'h98;
                    16'h3FD8: data_out = 8'h99;
                    16'h3FD9: data_out = 8'h9A;
                    16'h3FDA: data_out = 8'h9B;
                    16'h3FDB: data_out = 8'h9C;
                    16'h3FDC: data_out = 8'h9D;
                    16'h3FDD: data_out = 8'h9E;
                    16'h3FDE: data_out = 8'h9F;
                    16'h3FDF: data_out = 8'hA0;
                    16'h3FE0: data_out = 8'hA1;
                    16'h3FE1: data_out = 8'hA2;
                    16'h3FE2: data_out = 8'hA3;
                    16'h3FE3: data_out = 8'hA4;
                    16'h3FE4: data_out = 8'hA5;
                    16'h3FE5: data_out = 8'hA6;
                    16'h3FE6: data_out = 8'hA7;
                    16'h3FE7: data_out = 8'hA8;
                    16'h3FE8: data_out = 8'hA9;
                    16'h3FE9: data_out = 8'hAA;
                    16'h3FEA: data_out = 8'hAB;
                    16'h3FEB: data_out = 8'hAC;
                    16'h3FEC: data_out = 8'hAD;
                    16'h3FED: data_out = 8'hAE;
                    16'h3FEE: data_out = 8'hAF;
                    16'h3FEF: data_out = 8'hB0;
                    16'h3FF0: data_out = 8'hB1;
                    16'h3FF1: data_out = 8'hB2;
                    16'h3FF2: data_out = 8'hB3;
                    16'h3FF3: data_out = 8'hB4;
                    16'h3FF4: data_out = 8'hB5;
                    16'h3FF5: data_out = 8'hB6;
                    16'h3FF6: data_out = 8'hB7;
                    16'h3FF7: data_out = 8'hB8;
                    16'h3FF8: data_out = 8'hB9;
                    16'h3FF9: data_out = 8'hBA;
                    16'h3FFA: data_out = 8'hBB;
                    16'h3FFB: data_out = 8'hBC;
                    16'h3FFC: data_out = 8'hBD;
                    16'h3FFD: data_out = 8'hBE;
                    16'h3FFE: data_out = 8'hBF;
                    16'h3FFF: data_out = 8'hC0;
                    16'h4000: data_out = 8'h40;
                    16'h4001: data_out = 8'h41;
                    16'h4002: data_out = 8'h42;
                    16'h4003: data_out = 8'h43;
                    16'h4004: data_out = 8'h44;
                    16'h4005: data_out = 8'h45;
                    16'h4006: data_out = 8'h46;
                    16'h4007: data_out = 8'h47;
                    16'h4008: data_out = 8'h48;
                    16'h4009: data_out = 8'h49;
                    16'h400A: data_out = 8'h4A;
                    16'h400B: data_out = 8'h4B;
                    16'h400C: data_out = 8'h4C;
                    16'h400D: data_out = 8'h4D;
                    16'h400E: data_out = 8'h4E;
                    16'h400F: data_out = 8'h4F;
                    16'h4010: data_out = 8'h50;
                    16'h4011: data_out = 8'h51;
                    16'h4012: data_out = 8'h52;
                    16'h4013: data_out = 8'h53;
                    16'h4014: data_out = 8'h54;
                    16'h4015: data_out = 8'h55;
                    16'h4016: data_out = 8'h56;
                    16'h4017: data_out = 8'h57;
                    16'h4018: data_out = 8'h58;
                    16'h4019: data_out = 8'h59;
                    16'h401A: data_out = 8'h5A;
                    16'h401B: data_out = 8'h5B;
                    16'h401C: data_out = 8'h5C;
                    16'h401D: data_out = 8'h5D;
                    16'h401E: data_out = 8'h5E;
                    16'h401F: data_out = 8'h5F;
                    16'h4020: data_out = 8'h60;
                    16'h4021: data_out = 8'h61;
                    16'h4022: data_out = 8'h62;
                    16'h4023: data_out = 8'h63;
                    16'h4024: data_out = 8'h64;
                    16'h4025: data_out = 8'h65;
                    16'h4026: data_out = 8'h66;
                    16'h4027: data_out = 8'h67;
                    16'h4028: data_out = 8'h68;
                    16'h4029: data_out = 8'h69;
                    16'h402A: data_out = 8'h6A;
                    16'h402B: data_out = 8'h6B;
                    16'h402C: data_out = 8'h6C;
                    16'h402D: data_out = 8'h6D;
                    16'h402E: data_out = 8'h6E;
                    16'h402F: data_out = 8'h6F;
                    16'h4030: data_out = 8'h70;
                    16'h4031: data_out = 8'h71;
                    16'h4032: data_out = 8'h72;
                    16'h4033: data_out = 8'h73;
                    16'h4034: data_out = 8'h74;
                    16'h4035: data_out = 8'h75;
                    16'h4036: data_out = 8'h76;
                    16'h4037: data_out = 8'h77;
                    16'h4038: data_out = 8'h78;
                    16'h4039: data_out = 8'h79;
                    16'h403A: data_out = 8'h7A;
                    16'h403B: data_out = 8'h7B;
                    16'h403C: data_out = 8'h7C;
                    16'h403D: data_out = 8'h7D;
                    16'h403E: data_out = 8'h7E;
                    16'h403F: data_out = 8'h7F;
                    16'h4040: data_out = 8'h80;
                    16'h4041: data_out = 8'h81;
                    16'h4042: data_out = 8'h82;
                    16'h4043: data_out = 8'h83;
                    16'h4044: data_out = 8'h84;
                    16'h4045: data_out = 8'h85;
                    16'h4046: data_out = 8'h86;
                    16'h4047: data_out = 8'h87;
                    16'h4048: data_out = 8'h88;
                    16'h4049: data_out = 8'h89;
                    16'h404A: data_out = 8'h8A;
                    16'h404B: data_out = 8'h8B;
                    16'h404C: data_out = 8'h8C;
                    16'h404D: data_out = 8'h8D;
                    16'h404E: data_out = 8'h8E;
                    16'h404F: data_out = 8'h8F;
                    16'h4050: data_out = 8'h90;
                    16'h4051: data_out = 8'h91;
                    16'h4052: data_out = 8'h92;
                    16'h4053: data_out = 8'h93;
                    16'h4054: data_out = 8'h94;
                    16'h4055: data_out = 8'h95;
                    16'h4056: data_out = 8'h96;
                    16'h4057: data_out = 8'h97;
                    16'h4058: data_out = 8'h98;
                    16'h4059: data_out = 8'h99;
                    16'h405A: data_out = 8'h9A;
                    16'h405B: data_out = 8'h9B;
                    16'h405C: data_out = 8'h9C;
                    16'h405D: data_out = 8'h9D;
                    16'h405E: data_out = 8'h9E;
                    16'h405F: data_out = 8'h9F;
                    16'h4060: data_out = 8'hA0;
                    16'h4061: data_out = 8'hA1;
                    16'h4062: data_out = 8'hA2;
                    16'h4063: data_out = 8'hA3;
                    16'h4064: data_out = 8'hA4;
                    16'h4065: data_out = 8'hA5;
                    16'h4066: data_out = 8'hA6;
                    16'h4067: data_out = 8'hA7;
                    16'h4068: data_out = 8'hA8;
                    16'h4069: data_out = 8'hA9;
                    16'h406A: data_out = 8'hAA;
                    16'h406B: data_out = 8'hAB;
                    16'h406C: data_out = 8'hAC;
                    16'h406D: data_out = 8'hAD;
                    16'h406E: data_out = 8'hAE;
                    16'h406F: data_out = 8'hAF;
                    16'h4070: data_out = 8'hB0;
                    16'h4071: data_out = 8'hB1;
                    16'h4072: data_out = 8'hB2;
                    16'h4073: data_out = 8'hB3;
                    16'h4074: data_out = 8'hB4;
                    16'h4075: data_out = 8'hB5;
                    16'h4076: data_out = 8'hB6;
                    16'h4077: data_out = 8'hB7;
                    16'h4078: data_out = 8'hB8;
                    16'h4079: data_out = 8'hB9;
                    16'h407A: data_out = 8'hBA;
                    16'h407B: data_out = 8'hBB;
                    16'h407C: data_out = 8'hBC;
                    16'h407D: data_out = 8'hBD;
                    16'h407E: data_out = 8'hBE;
                    16'h407F: data_out = 8'hBF;
                    16'h4080: data_out = 8'h40;
                    16'h4081: data_out = 8'h3F;
                    16'h4082: data_out = 8'h3E;
                    16'h4083: data_out = 8'h3D;
                    16'h4084: data_out = 8'h3C;
                    16'h4085: data_out = 8'h3B;
                    16'h4086: data_out = 8'h3A;
                    16'h4087: data_out = 8'h39;
                    16'h4088: data_out = 8'h38;
                    16'h4089: data_out = 8'h37;
                    16'h408A: data_out = 8'h36;
                    16'h408B: data_out = 8'h35;
                    16'h408C: data_out = 8'h34;
                    16'h408D: data_out = 8'h33;
                    16'h408E: data_out = 8'h32;
                    16'h408F: data_out = 8'h31;
                    16'h4090: data_out = 8'h30;
                    16'h4091: data_out = 8'h2F;
                    16'h4092: data_out = 8'h2E;
                    16'h4093: data_out = 8'h2D;
                    16'h4094: data_out = 8'h2C;
                    16'h4095: data_out = 8'h2B;
                    16'h4096: data_out = 8'h2A;
                    16'h4097: data_out = 8'h29;
                    16'h4098: data_out = 8'h28;
                    16'h4099: data_out = 8'h27;
                    16'h409A: data_out = 8'h26;
                    16'h409B: data_out = 8'h25;
                    16'h409C: data_out = 8'h24;
                    16'h409D: data_out = 8'h23;
                    16'h409E: data_out = 8'h22;
                    16'h409F: data_out = 8'h21;
                    16'h40A0: data_out = 8'h20;
                    16'h40A1: data_out = 8'h1F;
                    16'h40A2: data_out = 8'h1E;
                    16'h40A3: data_out = 8'h1D;
                    16'h40A4: data_out = 8'h1C;
                    16'h40A5: data_out = 8'h1B;
                    16'h40A6: data_out = 8'h1A;
                    16'h40A7: data_out = 8'h19;
                    16'h40A8: data_out = 8'h18;
                    16'h40A9: data_out = 8'h17;
                    16'h40AA: data_out = 8'h16;
                    16'h40AB: data_out = 8'h15;
                    16'h40AC: data_out = 8'h14;
                    16'h40AD: data_out = 8'h13;
                    16'h40AE: data_out = 8'h12;
                    16'h40AF: data_out = 8'h11;
                    16'h40B0: data_out = 8'h10;
                    16'h40B1: data_out = 8'hF;
                    16'h40B2: data_out = 8'hE;
                    16'h40B3: data_out = 8'hD;
                    16'h40B4: data_out = 8'hC;
                    16'h40B5: data_out = 8'hB;
                    16'h40B6: data_out = 8'hA;
                    16'h40B7: data_out = 8'h9;
                    16'h40B8: data_out = 8'h8;
                    16'h40B9: data_out = 8'h7;
                    16'h40BA: data_out = 8'h6;
                    16'h40BB: data_out = 8'h5;
                    16'h40BC: data_out = 8'h4;
                    16'h40BD: data_out = 8'h3;
                    16'h40BE: data_out = 8'h2;
                    16'h40BF: data_out = 8'h1;
                    16'h40C0: data_out = 8'h0;
                    16'h40C1: data_out = 8'h81;
                    16'h40C2: data_out = 8'h82;
                    16'h40C3: data_out = 8'h83;
                    16'h40C4: data_out = 8'h84;
                    16'h40C5: data_out = 8'h85;
                    16'h40C6: data_out = 8'h86;
                    16'h40C7: data_out = 8'h87;
                    16'h40C8: data_out = 8'h88;
                    16'h40C9: data_out = 8'h89;
                    16'h40CA: data_out = 8'h8A;
                    16'h40CB: data_out = 8'h8B;
                    16'h40CC: data_out = 8'h8C;
                    16'h40CD: data_out = 8'h8D;
                    16'h40CE: data_out = 8'h8E;
                    16'h40CF: data_out = 8'h8F;
                    16'h40D0: data_out = 8'h90;
                    16'h40D1: data_out = 8'h91;
                    16'h40D2: data_out = 8'h92;
                    16'h40D3: data_out = 8'h93;
                    16'h40D4: data_out = 8'h94;
                    16'h40D5: data_out = 8'h95;
                    16'h40D6: data_out = 8'h96;
                    16'h40D7: data_out = 8'h97;
                    16'h40D8: data_out = 8'h98;
                    16'h40D9: data_out = 8'h99;
                    16'h40DA: data_out = 8'h9A;
                    16'h40DB: data_out = 8'h9B;
                    16'h40DC: data_out = 8'h9C;
                    16'h40DD: data_out = 8'h9D;
                    16'h40DE: data_out = 8'h9E;
                    16'h40DF: data_out = 8'h9F;
                    16'h40E0: data_out = 8'hA0;
                    16'h40E1: data_out = 8'hA1;
                    16'h40E2: data_out = 8'hA2;
                    16'h40E3: data_out = 8'hA3;
                    16'h40E4: data_out = 8'hA4;
                    16'h40E5: data_out = 8'hA5;
                    16'h40E6: data_out = 8'hA6;
                    16'h40E7: data_out = 8'hA7;
                    16'h40E8: data_out = 8'hA8;
                    16'h40E9: data_out = 8'hA9;
                    16'h40EA: data_out = 8'hAA;
                    16'h40EB: data_out = 8'hAB;
                    16'h40EC: data_out = 8'hAC;
                    16'h40ED: data_out = 8'hAD;
                    16'h40EE: data_out = 8'hAE;
                    16'h40EF: data_out = 8'hAF;
                    16'h40F0: data_out = 8'hB0;
                    16'h40F1: data_out = 8'hB1;
                    16'h40F2: data_out = 8'hB2;
                    16'h40F3: data_out = 8'hB3;
                    16'h40F4: data_out = 8'hB4;
                    16'h40F5: data_out = 8'hB5;
                    16'h40F6: data_out = 8'hB6;
                    16'h40F7: data_out = 8'hB7;
                    16'h40F8: data_out = 8'hB8;
                    16'h40F9: data_out = 8'hB9;
                    16'h40FA: data_out = 8'hBA;
                    16'h40FB: data_out = 8'hBB;
                    16'h40FC: data_out = 8'hBC;
                    16'h40FD: data_out = 8'hBD;
                    16'h40FE: data_out = 8'hBE;
                    16'h40FF: data_out = 8'hBF;
                    16'h4100: data_out = 8'h41;
                    16'h4101: data_out = 8'h42;
                    16'h4102: data_out = 8'h43;
                    16'h4103: data_out = 8'h44;
                    16'h4104: data_out = 8'h45;
                    16'h4105: data_out = 8'h46;
                    16'h4106: data_out = 8'h47;
                    16'h4107: data_out = 8'h48;
                    16'h4108: data_out = 8'h49;
                    16'h4109: data_out = 8'h4A;
                    16'h410A: data_out = 8'h4B;
                    16'h410B: data_out = 8'h4C;
                    16'h410C: data_out = 8'h4D;
                    16'h410D: data_out = 8'h4E;
                    16'h410E: data_out = 8'h4F;
                    16'h410F: data_out = 8'h50;
                    16'h4110: data_out = 8'h51;
                    16'h4111: data_out = 8'h52;
                    16'h4112: data_out = 8'h53;
                    16'h4113: data_out = 8'h54;
                    16'h4114: data_out = 8'h55;
                    16'h4115: data_out = 8'h56;
                    16'h4116: data_out = 8'h57;
                    16'h4117: data_out = 8'h58;
                    16'h4118: data_out = 8'h59;
                    16'h4119: data_out = 8'h5A;
                    16'h411A: data_out = 8'h5B;
                    16'h411B: data_out = 8'h5C;
                    16'h411C: data_out = 8'h5D;
                    16'h411D: data_out = 8'h5E;
                    16'h411E: data_out = 8'h5F;
                    16'h411F: data_out = 8'h60;
                    16'h4120: data_out = 8'h61;
                    16'h4121: data_out = 8'h62;
                    16'h4122: data_out = 8'h63;
                    16'h4123: data_out = 8'h64;
                    16'h4124: data_out = 8'h65;
                    16'h4125: data_out = 8'h66;
                    16'h4126: data_out = 8'h67;
                    16'h4127: data_out = 8'h68;
                    16'h4128: data_out = 8'h69;
                    16'h4129: data_out = 8'h6A;
                    16'h412A: data_out = 8'h6B;
                    16'h412B: data_out = 8'h6C;
                    16'h412C: data_out = 8'h6D;
                    16'h412D: data_out = 8'h6E;
                    16'h412E: data_out = 8'h6F;
                    16'h412F: data_out = 8'h70;
                    16'h4130: data_out = 8'h71;
                    16'h4131: data_out = 8'h72;
                    16'h4132: data_out = 8'h73;
                    16'h4133: data_out = 8'h74;
                    16'h4134: data_out = 8'h75;
                    16'h4135: data_out = 8'h76;
                    16'h4136: data_out = 8'h77;
                    16'h4137: data_out = 8'h78;
                    16'h4138: data_out = 8'h79;
                    16'h4139: data_out = 8'h7A;
                    16'h413A: data_out = 8'h7B;
                    16'h413B: data_out = 8'h7C;
                    16'h413C: data_out = 8'h7D;
                    16'h413D: data_out = 8'h7E;
                    16'h413E: data_out = 8'h7F;
                    16'h413F: data_out = 8'h80;
                    16'h4140: data_out = 8'h81;
                    16'h4141: data_out = 8'h82;
                    16'h4142: data_out = 8'h83;
                    16'h4143: data_out = 8'h84;
                    16'h4144: data_out = 8'h85;
                    16'h4145: data_out = 8'h86;
                    16'h4146: data_out = 8'h87;
                    16'h4147: data_out = 8'h88;
                    16'h4148: data_out = 8'h89;
                    16'h4149: data_out = 8'h8A;
                    16'h414A: data_out = 8'h8B;
                    16'h414B: data_out = 8'h8C;
                    16'h414C: data_out = 8'h8D;
                    16'h414D: data_out = 8'h8E;
                    16'h414E: data_out = 8'h8F;
                    16'h414F: data_out = 8'h90;
                    16'h4150: data_out = 8'h91;
                    16'h4151: data_out = 8'h92;
                    16'h4152: data_out = 8'h93;
                    16'h4153: data_out = 8'h94;
                    16'h4154: data_out = 8'h95;
                    16'h4155: data_out = 8'h96;
                    16'h4156: data_out = 8'h97;
                    16'h4157: data_out = 8'h98;
                    16'h4158: data_out = 8'h99;
                    16'h4159: data_out = 8'h9A;
                    16'h415A: data_out = 8'h9B;
                    16'h415B: data_out = 8'h9C;
                    16'h415C: data_out = 8'h9D;
                    16'h415D: data_out = 8'h9E;
                    16'h415E: data_out = 8'h9F;
                    16'h415F: data_out = 8'hA0;
                    16'h4160: data_out = 8'hA1;
                    16'h4161: data_out = 8'hA2;
                    16'h4162: data_out = 8'hA3;
                    16'h4163: data_out = 8'hA4;
                    16'h4164: data_out = 8'hA5;
                    16'h4165: data_out = 8'hA6;
                    16'h4166: data_out = 8'hA7;
                    16'h4167: data_out = 8'hA8;
                    16'h4168: data_out = 8'hA9;
                    16'h4169: data_out = 8'hAA;
                    16'h416A: data_out = 8'hAB;
                    16'h416B: data_out = 8'hAC;
                    16'h416C: data_out = 8'hAD;
                    16'h416D: data_out = 8'hAE;
                    16'h416E: data_out = 8'hAF;
                    16'h416F: data_out = 8'hB0;
                    16'h4170: data_out = 8'hB1;
                    16'h4171: data_out = 8'hB2;
                    16'h4172: data_out = 8'hB3;
                    16'h4173: data_out = 8'hB4;
                    16'h4174: data_out = 8'hB5;
                    16'h4175: data_out = 8'hB6;
                    16'h4176: data_out = 8'hB7;
                    16'h4177: data_out = 8'hB8;
                    16'h4178: data_out = 8'hB9;
                    16'h4179: data_out = 8'hBA;
                    16'h417A: data_out = 8'hBB;
                    16'h417B: data_out = 8'hBC;
                    16'h417C: data_out = 8'hBD;
                    16'h417D: data_out = 8'hBE;
                    16'h417E: data_out = 8'hBF;
                    16'h417F: data_out = 8'hC0;
                    16'h4180: data_out = 8'h41;
                    16'h4181: data_out = 8'h40;
                    16'h4182: data_out = 8'h3F;
                    16'h4183: data_out = 8'h3E;
                    16'h4184: data_out = 8'h3D;
                    16'h4185: data_out = 8'h3C;
                    16'h4186: data_out = 8'h3B;
                    16'h4187: data_out = 8'h3A;
                    16'h4188: data_out = 8'h39;
                    16'h4189: data_out = 8'h38;
                    16'h418A: data_out = 8'h37;
                    16'h418B: data_out = 8'h36;
                    16'h418C: data_out = 8'h35;
                    16'h418D: data_out = 8'h34;
                    16'h418E: data_out = 8'h33;
                    16'h418F: data_out = 8'h32;
                    16'h4190: data_out = 8'h31;
                    16'h4191: data_out = 8'h30;
                    16'h4192: data_out = 8'h2F;
                    16'h4193: data_out = 8'h2E;
                    16'h4194: data_out = 8'h2D;
                    16'h4195: data_out = 8'h2C;
                    16'h4196: data_out = 8'h2B;
                    16'h4197: data_out = 8'h2A;
                    16'h4198: data_out = 8'h29;
                    16'h4199: data_out = 8'h28;
                    16'h419A: data_out = 8'h27;
                    16'h419B: data_out = 8'h26;
                    16'h419C: data_out = 8'h25;
                    16'h419D: data_out = 8'h24;
                    16'h419E: data_out = 8'h23;
                    16'h419F: data_out = 8'h22;
                    16'h41A0: data_out = 8'h21;
                    16'h41A1: data_out = 8'h20;
                    16'h41A2: data_out = 8'h1F;
                    16'h41A3: data_out = 8'h1E;
                    16'h41A4: data_out = 8'h1D;
                    16'h41A5: data_out = 8'h1C;
                    16'h41A6: data_out = 8'h1B;
                    16'h41A7: data_out = 8'h1A;
                    16'h41A8: data_out = 8'h19;
                    16'h41A9: data_out = 8'h18;
                    16'h41AA: data_out = 8'h17;
                    16'h41AB: data_out = 8'h16;
                    16'h41AC: data_out = 8'h15;
                    16'h41AD: data_out = 8'h14;
                    16'h41AE: data_out = 8'h13;
                    16'h41AF: data_out = 8'h12;
                    16'h41B0: data_out = 8'h11;
                    16'h41B1: data_out = 8'h10;
                    16'h41B2: data_out = 8'hF;
                    16'h41B3: data_out = 8'hE;
                    16'h41B4: data_out = 8'hD;
                    16'h41B5: data_out = 8'hC;
                    16'h41B6: data_out = 8'hB;
                    16'h41B7: data_out = 8'hA;
                    16'h41B8: data_out = 8'h9;
                    16'h41B9: data_out = 8'h8;
                    16'h41BA: data_out = 8'h7;
                    16'h41BB: data_out = 8'h6;
                    16'h41BC: data_out = 8'h5;
                    16'h41BD: data_out = 8'h4;
                    16'h41BE: data_out = 8'h3;
                    16'h41BF: data_out = 8'h2;
                    16'h41C0: data_out = 8'h1;
                    16'h41C1: data_out = 8'h0;
                    16'h41C2: data_out = 8'h81;
                    16'h41C3: data_out = 8'h82;
                    16'h41C4: data_out = 8'h83;
                    16'h41C5: data_out = 8'h84;
                    16'h41C6: data_out = 8'h85;
                    16'h41C7: data_out = 8'h86;
                    16'h41C8: data_out = 8'h87;
                    16'h41C9: data_out = 8'h88;
                    16'h41CA: data_out = 8'h89;
                    16'h41CB: data_out = 8'h8A;
                    16'h41CC: data_out = 8'h8B;
                    16'h41CD: data_out = 8'h8C;
                    16'h41CE: data_out = 8'h8D;
                    16'h41CF: data_out = 8'h8E;
                    16'h41D0: data_out = 8'h8F;
                    16'h41D1: data_out = 8'h90;
                    16'h41D2: data_out = 8'h91;
                    16'h41D3: data_out = 8'h92;
                    16'h41D4: data_out = 8'h93;
                    16'h41D5: data_out = 8'h94;
                    16'h41D6: data_out = 8'h95;
                    16'h41D7: data_out = 8'h96;
                    16'h41D8: data_out = 8'h97;
                    16'h41D9: data_out = 8'h98;
                    16'h41DA: data_out = 8'h99;
                    16'h41DB: data_out = 8'h9A;
                    16'h41DC: data_out = 8'h9B;
                    16'h41DD: data_out = 8'h9C;
                    16'h41DE: data_out = 8'h9D;
                    16'h41DF: data_out = 8'h9E;
                    16'h41E0: data_out = 8'h9F;
                    16'h41E1: data_out = 8'hA0;
                    16'h41E2: data_out = 8'hA1;
                    16'h41E3: data_out = 8'hA2;
                    16'h41E4: data_out = 8'hA3;
                    16'h41E5: data_out = 8'hA4;
                    16'h41E6: data_out = 8'hA5;
                    16'h41E7: data_out = 8'hA6;
                    16'h41E8: data_out = 8'hA7;
                    16'h41E9: data_out = 8'hA8;
                    16'h41EA: data_out = 8'hA9;
                    16'h41EB: data_out = 8'hAA;
                    16'h41EC: data_out = 8'hAB;
                    16'h41ED: data_out = 8'hAC;
                    16'h41EE: data_out = 8'hAD;
                    16'h41EF: data_out = 8'hAE;
                    16'h41F0: data_out = 8'hAF;
                    16'h41F1: data_out = 8'hB0;
                    16'h41F2: data_out = 8'hB1;
                    16'h41F3: data_out = 8'hB2;
                    16'h41F4: data_out = 8'hB3;
                    16'h41F5: data_out = 8'hB4;
                    16'h41F6: data_out = 8'hB5;
                    16'h41F7: data_out = 8'hB6;
                    16'h41F8: data_out = 8'hB7;
                    16'h41F9: data_out = 8'hB8;
                    16'h41FA: data_out = 8'hB9;
                    16'h41FB: data_out = 8'hBA;
                    16'h41FC: data_out = 8'hBB;
                    16'h41FD: data_out = 8'hBC;
                    16'h41FE: data_out = 8'hBD;
                    16'h41FF: data_out = 8'hBE;
                    16'h4200: data_out = 8'h42;
                    16'h4201: data_out = 8'h43;
                    16'h4202: data_out = 8'h44;
                    16'h4203: data_out = 8'h45;
                    16'h4204: data_out = 8'h46;
                    16'h4205: data_out = 8'h47;
                    16'h4206: data_out = 8'h48;
                    16'h4207: data_out = 8'h49;
                    16'h4208: data_out = 8'h4A;
                    16'h4209: data_out = 8'h4B;
                    16'h420A: data_out = 8'h4C;
                    16'h420B: data_out = 8'h4D;
                    16'h420C: data_out = 8'h4E;
                    16'h420D: data_out = 8'h4F;
                    16'h420E: data_out = 8'h50;
                    16'h420F: data_out = 8'h51;
                    16'h4210: data_out = 8'h52;
                    16'h4211: data_out = 8'h53;
                    16'h4212: data_out = 8'h54;
                    16'h4213: data_out = 8'h55;
                    16'h4214: data_out = 8'h56;
                    16'h4215: data_out = 8'h57;
                    16'h4216: data_out = 8'h58;
                    16'h4217: data_out = 8'h59;
                    16'h4218: data_out = 8'h5A;
                    16'h4219: data_out = 8'h5B;
                    16'h421A: data_out = 8'h5C;
                    16'h421B: data_out = 8'h5D;
                    16'h421C: data_out = 8'h5E;
                    16'h421D: data_out = 8'h5F;
                    16'h421E: data_out = 8'h60;
                    16'h421F: data_out = 8'h61;
                    16'h4220: data_out = 8'h62;
                    16'h4221: data_out = 8'h63;
                    16'h4222: data_out = 8'h64;
                    16'h4223: data_out = 8'h65;
                    16'h4224: data_out = 8'h66;
                    16'h4225: data_out = 8'h67;
                    16'h4226: data_out = 8'h68;
                    16'h4227: data_out = 8'h69;
                    16'h4228: data_out = 8'h6A;
                    16'h4229: data_out = 8'h6B;
                    16'h422A: data_out = 8'h6C;
                    16'h422B: data_out = 8'h6D;
                    16'h422C: data_out = 8'h6E;
                    16'h422D: data_out = 8'h6F;
                    16'h422E: data_out = 8'h70;
                    16'h422F: data_out = 8'h71;
                    16'h4230: data_out = 8'h72;
                    16'h4231: data_out = 8'h73;
                    16'h4232: data_out = 8'h74;
                    16'h4233: data_out = 8'h75;
                    16'h4234: data_out = 8'h76;
                    16'h4235: data_out = 8'h77;
                    16'h4236: data_out = 8'h78;
                    16'h4237: data_out = 8'h79;
                    16'h4238: data_out = 8'h7A;
                    16'h4239: data_out = 8'h7B;
                    16'h423A: data_out = 8'h7C;
                    16'h423B: data_out = 8'h7D;
                    16'h423C: data_out = 8'h7E;
                    16'h423D: data_out = 8'h7F;
                    16'h423E: data_out = 8'h80;
                    16'h423F: data_out = 8'h81;
                    16'h4240: data_out = 8'h82;
                    16'h4241: data_out = 8'h83;
                    16'h4242: data_out = 8'h84;
                    16'h4243: data_out = 8'h85;
                    16'h4244: data_out = 8'h86;
                    16'h4245: data_out = 8'h87;
                    16'h4246: data_out = 8'h88;
                    16'h4247: data_out = 8'h89;
                    16'h4248: data_out = 8'h8A;
                    16'h4249: data_out = 8'h8B;
                    16'h424A: data_out = 8'h8C;
                    16'h424B: data_out = 8'h8D;
                    16'h424C: data_out = 8'h8E;
                    16'h424D: data_out = 8'h8F;
                    16'h424E: data_out = 8'h90;
                    16'h424F: data_out = 8'h91;
                    16'h4250: data_out = 8'h92;
                    16'h4251: data_out = 8'h93;
                    16'h4252: data_out = 8'h94;
                    16'h4253: data_out = 8'h95;
                    16'h4254: data_out = 8'h96;
                    16'h4255: data_out = 8'h97;
                    16'h4256: data_out = 8'h98;
                    16'h4257: data_out = 8'h99;
                    16'h4258: data_out = 8'h9A;
                    16'h4259: data_out = 8'h9B;
                    16'h425A: data_out = 8'h9C;
                    16'h425B: data_out = 8'h9D;
                    16'h425C: data_out = 8'h9E;
                    16'h425D: data_out = 8'h9F;
                    16'h425E: data_out = 8'hA0;
                    16'h425F: data_out = 8'hA1;
                    16'h4260: data_out = 8'hA2;
                    16'h4261: data_out = 8'hA3;
                    16'h4262: data_out = 8'hA4;
                    16'h4263: data_out = 8'hA5;
                    16'h4264: data_out = 8'hA6;
                    16'h4265: data_out = 8'hA7;
                    16'h4266: data_out = 8'hA8;
                    16'h4267: data_out = 8'hA9;
                    16'h4268: data_out = 8'hAA;
                    16'h4269: data_out = 8'hAB;
                    16'h426A: data_out = 8'hAC;
                    16'h426B: data_out = 8'hAD;
                    16'h426C: data_out = 8'hAE;
                    16'h426D: data_out = 8'hAF;
                    16'h426E: data_out = 8'hB0;
                    16'h426F: data_out = 8'hB1;
                    16'h4270: data_out = 8'hB2;
                    16'h4271: data_out = 8'hB3;
                    16'h4272: data_out = 8'hB4;
                    16'h4273: data_out = 8'hB5;
                    16'h4274: data_out = 8'hB6;
                    16'h4275: data_out = 8'hB7;
                    16'h4276: data_out = 8'hB8;
                    16'h4277: data_out = 8'hB9;
                    16'h4278: data_out = 8'hBA;
                    16'h4279: data_out = 8'hBB;
                    16'h427A: data_out = 8'hBC;
                    16'h427B: data_out = 8'hBD;
                    16'h427C: data_out = 8'hBE;
                    16'h427D: data_out = 8'hBF;
                    16'h427E: data_out = 8'hC0;
                    16'h427F: data_out = 8'hC1;
                    16'h4280: data_out = 8'h42;
                    16'h4281: data_out = 8'h41;
                    16'h4282: data_out = 8'h40;
                    16'h4283: data_out = 8'h3F;
                    16'h4284: data_out = 8'h3E;
                    16'h4285: data_out = 8'h3D;
                    16'h4286: data_out = 8'h3C;
                    16'h4287: data_out = 8'h3B;
                    16'h4288: data_out = 8'h3A;
                    16'h4289: data_out = 8'h39;
                    16'h428A: data_out = 8'h38;
                    16'h428B: data_out = 8'h37;
                    16'h428C: data_out = 8'h36;
                    16'h428D: data_out = 8'h35;
                    16'h428E: data_out = 8'h34;
                    16'h428F: data_out = 8'h33;
                    16'h4290: data_out = 8'h32;
                    16'h4291: data_out = 8'h31;
                    16'h4292: data_out = 8'h30;
                    16'h4293: data_out = 8'h2F;
                    16'h4294: data_out = 8'h2E;
                    16'h4295: data_out = 8'h2D;
                    16'h4296: data_out = 8'h2C;
                    16'h4297: data_out = 8'h2B;
                    16'h4298: data_out = 8'h2A;
                    16'h4299: data_out = 8'h29;
                    16'h429A: data_out = 8'h28;
                    16'h429B: data_out = 8'h27;
                    16'h429C: data_out = 8'h26;
                    16'h429D: data_out = 8'h25;
                    16'h429E: data_out = 8'h24;
                    16'h429F: data_out = 8'h23;
                    16'h42A0: data_out = 8'h22;
                    16'h42A1: data_out = 8'h21;
                    16'h42A2: data_out = 8'h20;
                    16'h42A3: data_out = 8'h1F;
                    16'h42A4: data_out = 8'h1E;
                    16'h42A5: data_out = 8'h1D;
                    16'h42A6: data_out = 8'h1C;
                    16'h42A7: data_out = 8'h1B;
                    16'h42A8: data_out = 8'h1A;
                    16'h42A9: data_out = 8'h19;
                    16'h42AA: data_out = 8'h18;
                    16'h42AB: data_out = 8'h17;
                    16'h42AC: data_out = 8'h16;
                    16'h42AD: data_out = 8'h15;
                    16'h42AE: data_out = 8'h14;
                    16'h42AF: data_out = 8'h13;
                    16'h42B0: data_out = 8'h12;
                    16'h42B1: data_out = 8'h11;
                    16'h42B2: data_out = 8'h10;
                    16'h42B3: data_out = 8'hF;
                    16'h42B4: data_out = 8'hE;
                    16'h42B5: data_out = 8'hD;
                    16'h42B6: data_out = 8'hC;
                    16'h42B7: data_out = 8'hB;
                    16'h42B8: data_out = 8'hA;
                    16'h42B9: data_out = 8'h9;
                    16'h42BA: data_out = 8'h8;
                    16'h42BB: data_out = 8'h7;
                    16'h42BC: data_out = 8'h6;
                    16'h42BD: data_out = 8'h5;
                    16'h42BE: data_out = 8'h4;
                    16'h42BF: data_out = 8'h3;
                    16'h42C0: data_out = 8'h2;
                    16'h42C1: data_out = 8'h1;
                    16'h42C2: data_out = 8'h0;
                    16'h42C3: data_out = 8'h81;
                    16'h42C4: data_out = 8'h82;
                    16'h42C5: data_out = 8'h83;
                    16'h42C6: data_out = 8'h84;
                    16'h42C7: data_out = 8'h85;
                    16'h42C8: data_out = 8'h86;
                    16'h42C9: data_out = 8'h87;
                    16'h42CA: data_out = 8'h88;
                    16'h42CB: data_out = 8'h89;
                    16'h42CC: data_out = 8'h8A;
                    16'h42CD: data_out = 8'h8B;
                    16'h42CE: data_out = 8'h8C;
                    16'h42CF: data_out = 8'h8D;
                    16'h42D0: data_out = 8'h8E;
                    16'h42D1: data_out = 8'h8F;
                    16'h42D2: data_out = 8'h90;
                    16'h42D3: data_out = 8'h91;
                    16'h42D4: data_out = 8'h92;
                    16'h42D5: data_out = 8'h93;
                    16'h42D6: data_out = 8'h94;
                    16'h42D7: data_out = 8'h95;
                    16'h42D8: data_out = 8'h96;
                    16'h42D9: data_out = 8'h97;
                    16'h42DA: data_out = 8'h98;
                    16'h42DB: data_out = 8'h99;
                    16'h42DC: data_out = 8'h9A;
                    16'h42DD: data_out = 8'h9B;
                    16'h42DE: data_out = 8'h9C;
                    16'h42DF: data_out = 8'h9D;
                    16'h42E0: data_out = 8'h9E;
                    16'h42E1: data_out = 8'h9F;
                    16'h42E2: data_out = 8'hA0;
                    16'h42E3: data_out = 8'hA1;
                    16'h42E4: data_out = 8'hA2;
                    16'h42E5: data_out = 8'hA3;
                    16'h42E6: data_out = 8'hA4;
                    16'h42E7: data_out = 8'hA5;
                    16'h42E8: data_out = 8'hA6;
                    16'h42E9: data_out = 8'hA7;
                    16'h42EA: data_out = 8'hA8;
                    16'h42EB: data_out = 8'hA9;
                    16'h42EC: data_out = 8'hAA;
                    16'h42ED: data_out = 8'hAB;
                    16'h42EE: data_out = 8'hAC;
                    16'h42EF: data_out = 8'hAD;
                    16'h42F0: data_out = 8'hAE;
                    16'h42F1: data_out = 8'hAF;
                    16'h42F2: data_out = 8'hB0;
                    16'h42F3: data_out = 8'hB1;
                    16'h42F4: data_out = 8'hB2;
                    16'h42F5: data_out = 8'hB3;
                    16'h42F6: data_out = 8'hB4;
                    16'h42F7: data_out = 8'hB5;
                    16'h42F8: data_out = 8'hB6;
                    16'h42F9: data_out = 8'hB7;
                    16'h42FA: data_out = 8'hB8;
                    16'h42FB: data_out = 8'hB9;
                    16'h42FC: data_out = 8'hBA;
                    16'h42FD: data_out = 8'hBB;
                    16'h42FE: data_out = 8'hBC;
                    16'h42FF: data_out = 8'hBD;
                    16'h4300: data_out = 8'h43;
                    16'h4301: data_out = 8'h44;
                    16'h4302: data_out = 8'h45;
                    16'h4303: data_out = 8'h46;
                    16'h4304: data_out = 8'h47;
                    16'h4305: data_out = 8'h48;
                    16'h4306: data_out = 8'h49;
                    16'h4307: data_out = 8'h4A;
                    16'h4308: data_out = 8'h4B;
                    16'h4309: data_out = 8'h4C;
                    16'h430A: data_out = 8'h4D;
                    16'h430B: data_out = 8'h4E;
                    16'h430C: data_out = 8'h4F;
                    16'h430D: data_out = 8'h50;
                    16'h430E: data_out = 8'h51;
                    16'h430F: data_out = 8'h52;
                    16'h4310: data_out = 8'h53;
                    16'h4311: data_out = 8'h54;
                    16'h4312: data_out = 8'h55;
                    16'h4313: data_out = 8'h56;
                    16'h4314: data_out = 8'h57;
                    16'h4315: data_out = 8'h58;
                    16'h4316: data_out = 8'h59;
                    16'h4317: data_out = 8'h5A;
                    16'h4318: data_out = 8'h5B;
                    16'h4319: data_out = 8'h5C;
                    16'h431A: data_out = 8'h5D;
                    16'h431B: data_out = 8'h5E;
                    16'h431C: data_out = 8'h5F;
                    16'h431D: data_out = 8'h60;
                    16'h431E: data_out = 8'h61;
                    16'h431F: data_out = 8'h62;
                    16'h4320: data_out = 8'h63;
                    16'h4321: data_out = 8'h64;
                    16'h4322: data_out = 8'h65;
                    16'h4323: data_out = 8'h66;
                    16'h4324: data_out = 8'h67;
                    16'h4325: data_out = 8'h68;
                    16'h4326: data_out = 8'h69;
                    16'h4327: data_out = 8'h6A;
                    16'h4328: data_out = 8'h6B;
                    16'h4329: data_out = 8'h6C;
                    16'h432A: data_out = 8'h6D;
                    16'h432B: data_out = 8'h6E;
                    16'h432C: data_out = 8'h6F;
                    16'h432D: data_out = 8'h70;
                    16'h432E: data_out = 8'h71;
                    16'h432F: data_out = 8'h72;
                    16'h4330: data_out = 8'h73;
                    16'h4331: data_out = 8'h74;
                    16'h4332: data_out = 8'h75;
                    16'h4333: data_out = 8'h76;
                    16'h4334: data_out = 8'h77;
                    16'h4335: data_out = 8'h78;
                    16'h4336: data_out = 8'h79;
                    16'h4337: data_out = 8'h7A;
                    16'h4338: data_out = 8'h7B;
                    16'h4339: data_out = 8'h7C;
                    16'h433A: data_out = 8'h7D;
                    16'h433B: data_out = 8'h7E;
                    16'h433C: data_out = 8'h7F;
                    16'h433D: data_out = 8'h80;
                    16'h433E: data_out = 8'h81;
                    16'h433F: data_out = 8'h82;
                    16'h4340: data_out = 8'h83;
                    16'h4341: data_out = 8'h84;
                    16'h4342: data_out = 8'h85;
                    16'h4343: data_out = 8'h86;
                    16'h4344: data_out = 8'h87;
                    16'h4345: data_out = 8'h88;
                    16'h4346: data_out = 8'h89;
                    16'h4347: data_out = 8'h8A;
                    16'h4348: data_out = 8'h8B;
                    16'h4349: data_out = 8'h8C;
                    16'h434A: data_out = 8'h8D;
                    16'h434B: data_out = 8'h8E;
                    16'h434C: data_out = 8'h8F;
                    16'h434D: data_out = 8'h90;
                    16'h434E: data_out = 8'h91;
                    16'h434F: data_out = 8'h92;
                    16'h4350: data_out = 8'h93;
                    16'h4351: data_out = 8'h94;
                    16'h4352: data_out = 8'h95;
                    16'h4353: data_out = 8'h96;
                    16'h4354: data_out = 8'h97;
                    16'h4355: data_out = 8'h98;
                    16'h4356: data_out = 8'h99;
                    16'h4357: data_out = 8'h9A;
                    16'h4358: data_out = 8'h9B;
                    16'h4359: data_out = 8'h9C;
                    16'h435A: data_out = 8'h9D;
                    16'h435B: data_out = 8'h9E;
                    16'h435C: data_out = 8'h9F;
                    16'h435D: data_out = 8'hA0;
                    16'h435E: data_out = 8'hA1;
                    16'h435F: data_out = 8'hA2;
                    16'h4360: data_out = 8'hA3;
                    16'h4361: data_out = 8'hA4;
                    16'h4362: data_out = 8'hA5;
                    16'h4363: data_out = 8'hA6;
                    16'h4364: data_out = 8'hA7;
                    16'h4365: data_out = 8'hA8;
                    16'h4366: data_out = 8'hA9;
                    16'h4367: data_out = 8'hAA;
                    16'h4368: data_out = 8'hAB;
                    16'h4369: data_out = 8'hAC;
                    16'h436A: data_out = 8'hAD;
                    16'h436B: data_out = 8'hAE;
                    16'h436C: data_out = 8'hAF;
                    16'h436D: data_out = 8'hB0;
                    16'h436E: data_out = 8'hB1;
                    16'h436F: data_out = 8'hB2;
                    16'h4370: data_out = 8'hB3;
                    16'h4371: data_out = 8'hB4;
                    16'h4372: data_out = 8'hB5;
                    16'h4373: data_out = 8'hB6;
                    16'h4374: data_out = 8'hB7;
                    16'h4375: data_out = 8'hB8;
                    16'h4376: data_out = 8'hB9;
                    16'h4377: data_out = 8'hBA;
                    16'h4378: data_out = 8'hBB;
                    16'h4379: data_out = 8'hBC;
                    16'h437A: data_out = 8'hBD;
                    16'h437B: data_out = 8'hBE;
                    16'h437C: data_out = 8'hBF;
                    16'h437D: data_out = 8'hC0;
                    16'h437E: data_out = 8'hC1;
                    16'h437F: data_out = 8'hC2;
                    16'h4380: data_out = 8'h43;
                    16'h4381: data_out = 8'h42;
                    16'h4382: data_out = 8'h41;
                    16'h4383: data_out = 8'h40;
                    16'h4384: data_out = 8'h3F;
                    16'h4385: data_out = 8'h3E;
                    16'h4386: data_out = 8'h3D;
                    16'h4387: data_out = 8'h3C;
                    16'h4388: data_out = 8'h3B;
                    16'h4389: data_out = 8'h3A;
                    16'h438A: data_out = 8'h39;
                    16'h438B: data_out = 8'h38;
                    16'h438C: data_out = 8'h37;
                    16'h438D: data_out = 8'h36;
                    16'h438E: data_out = 8'h35;
                    16'h438F: data_out = 8'h34;
                    16'h4390: data_out = 8'h33;
                    16'h4391: data_out = 8'h32;
                    16'h4392: data_out = 8'h31;
                    16'h4393: data_out = 8'h30;
                    16'h4394: data_out = 8'h2F;
                    16'h4395: data_out = 8'h2E;
                    16'h4396: data_out = 8'h2D;
                    16'h4397: data_out = 8'h2C;
                    16'h4398: data_out = 8'h2B;
                    16'h4399: data_out = 8'h2A;
                    16'h439A: data_out = 8'h29;
                    16'h439B: data_out = 8'h28;
                    16'h439C: data_out = 8'h27;
                    16'h439D: data_out = 8'h26;
                    16'h439E: data_out = 8'h25;
                    16'h439F: data_out = 8'h24;
                    16'h43A0: data_out = 8'h23;
                    16'h43A1: data_out = 8'h22;
                    16'h43A2: data_out = 8'h21;
                    16'h43A3: data_out = 8'h20;
                    16'h43A4: data_out = 8'h1F;
                    16'h43A5: data_out = 8'h1E;
                    16'h43A6: data_out = 8'h1D;
                    16'h43A7: data_out = 8'h1C;
                    16'h43A8: data_out = 8'h1B;
                    16'h43A9: data_out = 8'h1A;
                    16'h43AA: data_out = 8'h19;
                    16'h43AB: data_out = 8'h18;
                    16'h43AC: data_out = 8'h17;
                    16'h43AD: data_out = 8'h16;
                    16'h43AE: data_out = 8'h15;
                    16'h43AF: data_out = 8'h14;
                    16'h43B0: data_out = 8'h13;
                    16'h43B1: data_out = 8'h12;
                    16'h43B2: data_out = 8'h11;
                    16'h43B3: data_out = 8'h10;
                    16'h43B4: data_out = 8'hF;
                    16'h43B5: data_out = 8'hE;
                    16'h43B6: data_out = 8'hD;
                    16'h43B7: data_out = 8'hC;
                    16'h43B8: data_out = 8'hB;
                    16'h43B9: data_out = 8'hA;
                    16'h43BA: data_out = 8'h9;
                    16'h43BB: data_out = 8'h8;
                    16'h43BC: data_out = 8'h7;
                    16'h43BD: data_out = 8'h6;
                    16'h43BE: data_out = 8'h5;
                    16'h43BF: data_out = 8'h4;
                    16'h43C0: data_out = 8'h3;
                    16'h43C1: data_out = 8'h2;
                    16'h43C2: data_out = 8'h1;
                    16'h43C3: data_out = 8'h0;
                    16'h43C4: data_out = 8'h81;
                    16'h43C5: data_out = 8'h82;
                    16'h43C6: data_out = 8'h83;
                    16'h43C7: data_out = 8'h84;
                    16'h43C8: data_out = 8'h85;
                    16'h43C9: data_out = 8'h86;
                    16'h43CA: data_out = 8'h87;
                    16'h43CB: data_out = 8'h88;
                    16'h43CC: data_out = 8'h89;
                    16'h43CD: data_out = 8'h8A;
                    16'h43CE: data_out = 8'h8B;
                    16'h43CF: data_out = 8'h8C;
                    16'h43D0: data_out = 8'h8D;
                    16'h43D1: data_out = 8'h8E;
                    16'h43D2: data_out = 8'h8F;
                    16'h43D3: data_out = 8'h90;
                    16'h43D4: data_out = 8'h91;
                    16'h43D5: data_out = 8'h92;
                    16'h43D6: data_out = 8'h93;
                    16'h43D7: data_out = 8'h94;
                    16'h43D8: data_out = 8'h95;
                    16'h43D9: data_out = 8'h96;
                    16'h43DA: data_out = 8'h97;
                    16'h43DB: data_out = 8'h98;
                    16'h43DC: data_out = 8'h99;
                    16'h43DD: data_out = 8'h9A;
                    16'h43DE: data_out = 8'h9B;
                    16'h43DF: data_out = 8'h9C;
                    16'h43E0: data_out = 8'h9D;
                    16'h43E1: data_out = 8'h9E;
                    16'h43E2: data_out = 8'h9F;
                    16'h43E3: data_out = 8'hA0;
                    16'h43E4: data_out = 8'hA1;
                    16'h43E5: data_out = 8'hA2;
                    16'h43E6: data_out = 8'hA3;
                    16'h43E7: data_out = 8'hA4;
                    16'h43E8: data_out = 8'hA5;
                    16'h43E9: data_out = 8'hA6;
                    16'h43EA: data_out = 8'hA7;
                    16'h43EB: data_out = 8'hA8;
                    16'h43EC: data_out = 8'hA9;
                    16'h43ED: data_out = 8'hAA;
                    16'h43EE: data_out = 8'hAB;
                    16'h43EF: data_out = 8'hAC;
                    16'h43F0: data_out = 8'hAD;
                    16'h43F1: data_out = 8'hAE;
                    16'h43F2: data_out = 8'hAF;
                    16'h43F3: data_out = 8'hB0;
                    16'h43F4: data_out = 8'hB1;
                    16'h43F5: data_out = 8'hB2;
                    16'h43F6: data_out = 8'hB3;
                    16'h43F7: data_out = 8'hB4;
                    16'h43F8: data_out = 8'hB5;
                    16'h43F9: data_out = 8'hB6;
                    16'h43FA: data_out = 8'hB7;
                    16'h43FB: data_out = 8'hB8;
                    16'h43FC: data_out = 8'hB9;
                    16'h43FD: data_out = 8'hBA;
                    16'h43FE: data_out = 8'hBB;
                    16'h43FF: data_out = 8'hBC;
                    16'h4400: data_out = 8'h44;
                    16'h4401: data_out = 8'h45;
                    16'h4402: data_out = 8'h46;
                    16'h4403: data_out = 8'h47;
                    16'h4404: data_out = 8'h48;
                    16'h4405: data_out = 8'h49;
                    16'h4406: data_out = 8'h4A;
                    16'h4407: data_out = 8'h4B;
                    16'h4408: data_out = 8'h4C;
                    16'h4409: data_out = 8'h4D;
                    16'h440A: data_out = 8'h4E;
                    16'h440B: data_out = 8'h4F;
                    16'h440C: data_out = 8'h50;
                    16'h440D: data_out = 8'h51;
                    16'h440E: data_out = 8'h52;
                    16'h440F: data_out = 8'h53;
                    16'h4410: data_out = 8'h54;
                    16'h4411: data_out = 8'h55;
                    16'h4412: data_out = 8'h56;
                    16'h4413: data_out = 8'h57;
                    16'h4414: data_out = 8'h58;
                    16'h4415: data_out = 8'h59;
                    16'h4416: data_out = 8'h5A;
                    16'h4417: data_out = 8'h5B;
                    16'h4418: data_out = 8'h5C;
                    16'h4419: data_out = 8'h5D;
                    16'h441A: data_out = 8'h5E;
                    16'h441B: data_out = 8'h5F;
                    16'h441C: data_out = 8'h60;
                    16'h441D: data_out = 8'h61;
                    16'h441E: data_out = 8'h62;
                    16'h441F: data_out = 8'h63;
                    16'h4420: data_out = 8'h64;
                    16'h4421: data_out = 8'h65;
                    16'h4422: data_out = 8'h66;
                    16'h4423: data_out = 8'h67;
                    16'h4424: data_out = 8'h68;
                    16'h4425: data_out = 8'h69;
                    16'h4426: data_out = 8'h6A;
                    16'h4427: data_out = 8'h6B;
                    16'h4428: data_out = 8'h6C;
                    16'h4429: data_out = 8'h6D;
                    16'h442A: data_out = 8'h6E;
                    16'h442B: data_out = 8'h6F;
                    16'h442C: data_out = 8'h70;
                    16'h442D: data_out = 8'h71;
                    16'h442E: data_out = 8'h72;
                    16'h442F: data_out = 8'h73;
                    16'h4430: data_out = 8'h74;
                    16'h4431: data_out = 8'h75;
                    16'h4432: data_out = 8'h76;
                    16'h4433: data_out = 8'h77;
                    16'h4434: data_out = 8'h78;
                    16'h4435: data_out = 8'h79;
                    16'h4436: data_out = 8'h7A;
                    16'h4437: data_out = 8'h7B;
                    16'h4438: data_out = 8'h7C;
                    16'h4439: data_out = 8'h7D;
                    16'h443A: data_out = 8'h7E;
                    16'h443B: data_out = 8'h7F;
                    16'h443C: data_out = 8'h80;
                    16'h443D: data_out = 8'h81;
                    16'h443E: data_out = 8'h82;
                    16'h443F: data_out = 8'h83;
                    16'h4440: data_out = 8'h84;
                    16'h4441: data_out = 8'h85;
                    16'h4442: data_out = 8'h86;
                    16'h4443: data_out = 8'h87;
                    16'h4444: data_out = 8'h88;
                    16'h4445: data_out = 8'h89;
                    16'h4446: data_out = 8'h8A;
                    16'h4447: data_out = 8'h8B;
                    16'h4448: data_out = 8'h8C;
                    16'h4449: data_out = 8'h8D;
                    16'h444A: data_out = 8'h8E;
                    16'h444B: data_out = 8'h8F;
                    16'h444C: data_out = 8'h90;
                    16'h444D: data_out = 8'h91;
                    16'h444E: data_out = 8'h92;
                    16'h444F: data_out = 8'h93;
                    16'h4450: data_out = 8'h94;
                    16'h4451: data_out = 8'h95;
                    16'h4452: data_out = 8'h96;
                    16'h4453: data_out = 8'h97;
                    16'h4454: data_out = 8'h98;
                    16'h4455: data_out = 8'h99;
                    16'h4456: data_out = 8'h9A;
                    16'h4457: data_out = 8'h9B;
                    16'h4458: data_out = 8'h9C;
                    16'h4459: data_out = 8'h9D;
                    16'h445A: data_out = 8'h9E;
                    16'h445B: data_out = 8'h9F;
                    16'h445C: data_out = 8'hA0;
                    16'h445D: data_out = 8'hA1;
                    16'h445E: data_out = 8'hA2;
                    16'h445F: data_out = 8'hA3;
                    16'h4460: data_out = 8'hA4;
                    16'h4461: data_out = 8'hA5;
                    16'h4462: data_out = 8'hA6;
                    16'h4463: data_out = 8'hA7;
                    16'h4464: data_out = 8'hA8;
                    16'h4465: data_out = 8'hA9;
                    16'h4466: data_out = 8'hAA;
                    16'h4467: data_out = 8'hAB;
                    16'h4468: data_out = 8'hAC;
                    16'h4469: data_out = 8'hAD;
                    16'h446A: data_out = 8'hAE;
                    16'h446B: data_out = 8'hAF;
                    16'h446C: data_out = 8'hB0;
                    16'h446D: data_out = 8'hB1;
                    16'h446E: data_out = 8'hB2;
                    16'h446F: data_out = 8'hB3;
                    16'h4470: data_out = 8'hB4;
                    16'h4471: data_out = 8'hB5;
                    16'h4472: data_out = 8'hB6;
                    16'h4473: data_out = 8'hB7;
                    16'h4474: data_out = 8'hB8;
                    16'h4475: data_out = 8'hB9;
                    16'h4476: data_out = 8'hBA;
                    16'h4477: data_out = 8'hBB;
                    16'h4478: data_out = 8'hBC;
                    16'h4479: data_out = 8'hBD;
                    16'h447A: data_out = 8'hBE;
                    16'h447B: data_out = 8'hBF;
                    16'h447C: data_out = 8'hC0;
                    16'h447D: data_out = 8'hC1;
                    16'h447E: data_out = 8'hC2;
                    16'h447F: data_out = 8'hC3;
                    16'h4480: data_out = 8'h44;
                    16'h4481: data_out = 8'h43;
                    16'h4482: data_out = 8'h42;
                    16'h4483: data_out = 8'h41;
                    16'h4484: data_out = 8'h40;
                    16'h4485: data_out = 8'h3F;
                    16'h4486: data_out = 8'h3E;
                    16'h4487: data_out = 8'h3D;
                    16'h4488: data_out = 8'h3C;
                    16'h4489: data_out = 8'h3B;
                    16'h448A: data_out = 8'h3A;
                    16'h448B: data_out = 8'h39;
                    16'h448C: data_out = 8'h38;
                    16'h448D: data_out = 8'h37;
                    16'h448E: data_out = 8'h36;
                    16'h448F: data_out = 8'h35;
                    16'h4490: data_out = 8'h34;
                    16'h4491: data_out = 8'h33;
                    16'h4492: data_out = 8'h32;
                    16'h4493: data_out = 8'h31;
                    16'h4494: data_out = 8'h30;
                    16'h4495: data_out = 8'h2F;
                    16'h4496: data_out = 8'h2E;
                    16'h4497: data_out = 8'h2D;
                    16'h4498: data_out = 8'h2C;
                    16'h4499: data_out = 8'h2B;
                    16'h449A: data_out = 8'h2A;
                    16'h449B: data_out = 8'h29;
                    16'h449C: data_out = 8'h28;
                    16'h449D: data_out = 8'h27;
                    16'h449E: data_out = 8'h26;
                    16'h449F: data_out = 8'h25;
                    16'h44A0: data_out = 8'h24;
                    16'h44A1: data_out = 8'h23;
                    16'h44A2: data_out = 8'h22;
                    16'h44A3: data_out = 8'h21;
                    16'h44A4: data_out = 8'h20;
                    16'h44A5: data_out = 8'h1F;
                    16'h44A6: data_out = 8'h1E;
                    16'h44A7: data_out = 8'h1D;
                    16'h44A8: data_out = 8'h1C;
                    16'h44A9: data_out = 8'h1B;
                    16'h44AA: data_out = 8'h1A;
                    16'h44AB: data_out = 8'h19;
                    16'h44AC: data_out = 8'h18;
                    16'h44AD: data_out = 8'h17;
                    16'h44AE: data_out = 8'h16;
                    16'h44AF: data_out = 8'h15;
                    16'h44B0: data_out = 8'h14;
                    16'h44B1: data_out = 8'h13;
                    16'h44B2: data_out = 8'h12;
                    16'h44B3: data_out = 8'h11;
                    16'h44B4: data_out = 8'h10;
                    16'h44B5: data_out = 8'hF;
                    16'h44B6: data_out = 8'hE;
                    16'h44B7: data_out = 8'hD;
                    16'h44B8: data_out = 8'hC;
                    16'h44B9: data_out = 8'hB;
                    16'h44BA: data_out = 8'hA;
                    16'h44BB: data_out = 8'h9;
                    16'h44BC: data_out = 8'h8;
                    16'h44BD: data_out = 8'h7;
                    16'h44BE: data_out = 8'h6;
                    16'h44BF: data_out = 8'h5;
                    16'h44C0: data_out = 8'h4;
                    16'h44C1: data_out = 8'h3;
                    16'h44C2: data_out = 8'h2;
                    16'h44C3: data_out = 8'h1;
                    16'h44C4: data_out = 8'h0;
                    16'h44C5: data_out = 8'h81;
                    16'h44C6: data_out = 8'h82;
                    16'h44C7: data_out = 8'h83;
                    16'h44C8: data_out = 8'h84;
                    16'h44C9: data_out = 8'h85;
                    16'h44CA: data_out = 8'h86;
                    16'h44CB: data_out = 8'h87;
                    16'h44CC: data_out = 8'h88;
                    16'h44CD: data_out = 8'h89;
                    16'h44CE: data_out = 8'h8A;
                    16'h44CF: data_out = 8'h8B;
                    16'h44D0: data_out = 8'h8C;
                    16'h44D1: data_out = 8'h8D;
                    16'h44D2: data_out = 8'h8E;
                    16'h44D3: data_out = 8'h8F;
                    16'h44D4: data_out = 8'h90;
                    16'h44D5: data_out = 8'h91;
                    16'h44D6: data_out = 8'h92;
                    16'h44D7: data_out = 8'h93;
                    16'h44D8: data_out = 8'h94;
                    16'h44D9: data_out = 8'h95;
                    16'h44DA: data_out = 8'h96;
                    16'h44DB: data_out = 8'h97;
                    16'h44DC: data_out = 8'h98;
                    16'h44DD: data_out = 8'h99;
                    16'h44DE: data_out = 8'h9A;
                    16'h44DF: data_out = 8'h9B;
                    16'h44E0: data_out = 8'h9C;
                    16'h44E1: data_out = 8'h9D;
                    16'h44E2: data_out = 8'h9E;
                    16'h44E3: data_out = 8'h9F;
                    16'h44E4: data_out = 8'hA0;
                    16'h44E5: data_out = 8'hA1;
                    16'h44E6: data_out = 8'hA2;
                    16'h44E7: data_out = 8'hA3;
                    16'h44E8: data_out = 8'hA4;
                    16'h44E9: data_out = 8'hA5;
                    16'h44EA: data_out = 8'hA6;
                    16'h44EB: data_out = 8'hA7;
                    16'h44EC: data_out = 8'hA8;
                    16'h44ED: data_out = 8'hA9;
                    16'h44EE: data_out = 8'hAA;
                    16'h44EF: data_out = 8'hAB;
                    16'h44F0: data_out = 8'hAC;
                    16'h44F1: data_out = 8'hAD;
                    16'h44F2: data_out = 8'hAE;
                    16'h44F3: data_out = 8'hAF;
                    16'h44F4: data_out = 8'hB0;
                    16'h44F5: data_out = 8'hB1;
                    16'h44F6: data_out = 8'hB2;
                    16'h44F7: data_out = 8'hB3;
                    16'h44F8: data_out = 8'hB4;
                    16'h44F9: data_out = 8'hB5;
                    16'h44FA: data_out = 8'hB6;
                    16'h44FB: data_out = 8'hB7;
                    16'h44FC: data_out = 8'hB8;
                    16'h44FD: data_out = 8'hB9;
                    16'h44FE: data_out = 8'hBA;
                    16'h44FF: data_out = 8'hBB;
                    16'h4500: data_out = 8'h45;
                    16'h4501: data_out = 8'h46;
                    16'h4502: data_out = 8'h47;
                    16'h4503: data_out = 8'h48;
                    16'h4504: data_out = 8'h49;
                    16'h4505: data_out = 8'h4A;
                    16'h4506: data_out = 8'h4B;
                    16'h4507: data_out = 8'h4C;
                    16'h4508: data_out = 8'h4D;
                    16'h4509: data_out = 8'h4E;
                    16'h450A: data_out = 8'h4F;
                    16'h450B: data_out = 8'h50;
                    16'h450C: data_out = 8'h51;
                    16'h450D: data_out = 8'h52;
                    16'h450E: data_out = 8'h53;
                    16'h450F: data_out = 8'h54;
                    16'h4510: data_out = 8'h55;
                    16'h4511: data_out = 8'h56;
                    16'h4512: data_out = 8'h57;
                    16'h4513: data_out = 8'h58;
                    16'h4514: data_out = 8'h59;
                    16'h4515: data_out = 8'h5A;
                    16'h4516: data_out = 8'h5B;
                    16'h4517: data_out = 8'h5C;
                    16'h4518: data_out = 8'h5D;
                    16'h4519: data_out = 8'h5E;
                    16'h451A: data_out = 8'h5F;
                    16'h451B: data_out = 8'h60;
                    16'h451C: data_out = 8'h61;
                    16'h451D: data_out = 8'h62;
                    16'h451E: data_out = 8'h63;
                    16'h451F: data_out = 8'h64;
                    16'h4520: data_out = 8'h65;
                    16'h4521: data_out = 8'h66;
                    16'h4522: data_out = 8'h67;
                    16'h4523: data_out = 8'h68;
                    16'h4524: data_out = 8'h69;
                    16'h4525: data_out = 8'h6A;
                    16'h4526: data_out = 8'h6B;
                    16'h4527: data_out = 8'h6C;
                    16'h4528: data_out = 8'h6D;
                    16'h4529: data_out = 8'h6E;
                    16'h452A: data_out = 8'h6F;
                    16'h452B: data_out = 8'h70;
                    16'h452C: data_out = 8'h71;
                    16'h452D: data_out = 8'h72;
                    16'h452E: data_out = 8'h73;
                    16'h452F: data_out = 8'h74;
                    16'h4530: data_out = 8'h75;
                    16'h4531: data_out = 8'h76;
                    16'h4532: data_out = 8'h77;
                    16'h4533: data_out = 8'h78;
                    16'h4534: data_out = 8'h79;
                    16'h4535: data_out = 8'h7A;
                    16'h4536: data_out = 8'h7B;
                    16'h4537: data_out = 8'h7C;
                    16'h4538: data_out = 8'h7D;
                    16'h4539: data_out = 8'h7E;
                    16'h453A: data_out = 8'h7F;
                    16'h453B: data_out = 8'h80;
                    16'h453C: data_out = 8'h81;
                    16'h453D: data_out = 8'h82;
                    16'h453E: data_out = 8'h83;
                    16'h453F: data_out = 8'h84;
                    16'h4540: data_out = 8'h85;
                    16'h4541: data_out = 8'h86;
                    16'h4542: data_out = 8'h87;
                    16'h4543: data_out = 8'h88;
                    16'h4544: data_out = 8'h89;
                    16'h4545: data_out = 8'h8A;
                    16'h4546: data_out = 8'h8B;
                    16'h4547: data_out = 8'h8C;
                    16'h4548: data_out = 8'h8D;
                    16'h4549: data_out = 8'h8E;
                    16'h454A: data_out = 8'h8F;
                    16'h454B: data_out = 8'h90;
                    16'h454C: data_out = 8'h91;
                    16'h454D: data_out = 8'h92;
                    16'h454E: data_out = 8'h93;
                    16'h454F: data_out = 8'h94;
                    16'h4550: data_out = 8'h95;
                    16'h4551: data_out = 8'h96;
                    16'h4552: data_out = 8'h97;
                    16'h4553: data_out = 8'h98;
                    16'h4554: data_out = 8'h99;
                    16'h4555: data_out = 8'h9A;
                    16'h4556: data_out = 8'h9B;
                    16'h4557: data_out = 8'h9C;
                    16'h4558: data_out = 8'h9D;
                    16'h4559: data_out = 8'h9E;
                    16'h455A: data_out = 8'h9F;
                    16'h455B: data_out = 8'hA0;
                    16'h455C: data_out = 8'hA1;
                    16'h455D: data_out = 8'hA2;
                    16'h455E: data_out = 8'hA3;
                    16'h455F: data_out = 8'hA4;
                    16'h4560: data_out = 8'hA5;
                    16'h4561: data_out = 8'hA6;
                    16'h4562: data_out = 8'hA7;
                    16'h4563: data_out = 8'hA8;
                    16'h4564: data_out = 8'hA9;
                    16'h4565: data_out = 8'hAA;
                    16'h4566: data_out = 8'hAB;
                    16'h4567: data_out = 8'hAC;
                    16'h4568: data_out = 8'hAD;
                    16'h4569: data_out = 8'hAE;
                    16'h456A: data_out = 8'hAF;
                    16'h456B: data_out = 8'hB0;
                    16'h456C: data_out = 8'hB1;
                    16'h456D: data_out = 8'hB2;
                    16'h456E: data_out = 8'hB3;
                    16'h456F: data_out = 8'hB4;
                    16'h4570: data_out = 8'hB5;
                    16'h4571: data_out = 8'hB6;
                    16'h4572: data_out = 8'hB7;
                    16'h4573: data_out = 8'hB8;
                    16'h4574: data_out = 8'hB9;
                    16'h4575: data_out = 8'hBA;
                    16'h4576: data_out = 8'hBB;
                    16'h4577: data_out = 8'hBC;
                    16'h4578: data_out = 8'hBD;
                    16'h4579: data_out = 8'hBE;
                    16'h457A: data_out = 8'hBF;
                    16'h457B: data_out = 8'hC0;
                    16'h457C: data_out = 8'hC1;
                    16'h457D: data_out = 8'hC2;
                    16'h457E: data_out = 8'hC3;
                    16'h457F: data_out = 8'hC4;
                    16'h4580: data_out = 8'h45;
                    16'h4581: data_out = 8'h44;
                    16'h4582: data_out = 8'h43;
                    16'h4583: data_out = 8'h42;
                    16'h4584: data_out = 8'h41;
                    16'h4585: data_out = 8'h40;
                    16'h4586: data_out = 8'h3F;
                    16'h4587: data_out = 8'h3E;
                    16'h4588: data_out = 8'h3D;
                    16'h4589: data_out = 8'h3C;
                    16'h458A: data_out = 8'h3B;
                    16'h458B: data_out = 8'h3A;
                    16'h458C: data_out = 8'h39;
                    16'h458D: data_out = 8'h38;
                    16'h458E: data_out = 8'h37;
                    16'h458F: data_out = 8'h36;
                    16'h4590: data_out = 8'h35;
                    16'h4591: data_out = 8'h34;
                    16'h4592: data_out = 8'h33;
                    16'h4593: data_out = 8'h32;
                    16'h4594: data_out = 8'h31;
                    16'h4595: data_out = 8'h30;
                    16'h4596: data_out = 8'h2F;
                    16'h4597: data_out = 8'h2E;
                    16'h4598: data_out = 8'h2D;
                    16'h4599: data_out = 8'h2C;
                    16'h459A: data_out = 8'h2B;
                    16'h459B: data_out = 8'h2A;
                    16'h459C: data_out = 8'h29;
                    16'h459D: data_out = 8'h28;
                    16'h459E: data_out = 8'h27;
                    16'h459F: data_out = 8'h26;
                    16'h45A0: data_out = 8'h25;
                    16'h45A1: data_out = 8'h24;
                    16'h45A2: data_out = 8'h23;
                    16'h45A3: data_out = 8'h22;
                    16'h45A4: data_out = 8'h21;
                    16'h45A5: data_out = 8'h20;
                    16'h45A6: data_out = 8'h1F;
                    16'h45A7: data_out = 8'h1E;
                    16'h45A8: data_out = 8'h1D;
                    16'h45A9: data_out = 8'h1C;
                    16'h45AA: data_out = 8'h1B;
                    16'h45AB: data_out = 8'h1A;
                    16'h45AC: data_out = 8'h19;
                    16'h45AD: data_out = 8'h18;
                    16'h45AE: data_out = 8'h17;
                    16'h45AF: data_out = 8'h16;
                    16'h45B0: data_out = 8'h15;
                    16'h45B1: data_out = 8'h14;
                    16'h45B2: data_out = 8'h13;
                    16'h45B3: data_out = 8'h12;
                    16'h45B4: data_out = 8'h11;
                    16'h45B5: data_out = 8'h10;
                    16'h45B6: data_out = 8'hF;
                    16'h45B7: data_out = 8'hE;
                    16'h45B8: data_out = 8'hD;
                    16'h45B9: data_out = 8'hC;
                    16'h45BA: data_out = 8'hB;
                    16'h45BB: data_out = 8'hA;
                    16'h45BC: data_out = 8'h9;
                    16'h45BD: data_out = 8'h8;
                    16'h45BE: data_out = 8'h7;
                    16'h45BF: data_out = 8'h6;
                    16'h45C0: data_out = 8'h5;
                    16'h45C1: data_out = 8'h4;
                    16'h45C2: data_out = 8'h3;
                    16'h45C3: data_out = 8'h2;
                    16'h45C4: data_out = 8'h1;
                    16'h45C5: data_out = 8'h0;
                    16'h45C6: data_out = 8'h81;
                    16'h45C7: data_out = 8'h82;
                    16'h45C8: data_out = 8'h83;
                    16'h45C9: data_out = 8'h84;
                    16'h45CA: data_out = 8'h85;
                    16'h45CB: data_out = 8'h86;
                    16'h45CC: data_out = 8'h87;
                    16'h45CD: data_out = 8'h88;
                    16'h45CE: data_out = 8'h89;
                    16'h45CF: data_out = 8'h8A;
                    16'h45D0: data_out = 8'h8B;
                    16'h45D1: data_out = 8'h8C;
                    16'h45D2: data_out = 8'h8D;
                    16'h45D3: data_out = 8'h8E;
                    16'h45D4: data_out = 8'h8F;
                    16'h45D5: data_out = 8'h90;
                    16'h45D6: data_out = 8'h91;
                    16'h45D7: data_out = 8'h92;
                    16'h45D8: data_out = 8'h93;
                    16'h45D9: data_out = 8'h94;
                    16'h45DA: data_out = 8'h95;
                    16'h45DB: data_out = 8'h96;
                    16'h45DC: data_out = 8'h97;
                    16'h45DD: data_out = 8'h98;
                    16'h45DE: data_out = 8'h99;
                    16'h45DF: data_out = 8'h9A;
                    16'h45E0: data_out = 8'h9B;
                    16'h45E1: data_out = 8'h9C;
                    16'h45E2: data_out = 8'h9D;
                    16'h45E3: data_out = 8'h9E;
                    16'h45E4: data_out = 8'h9F;
                    16'h45E5: data_out = 8'hA0;
                    16'h45E6: data_out = 8'hA1;
                    16'h45E7: data_out = 8'hA2;
                    16'h45E8: data_out = 8'hA3;
                    16'h45E9: data_out = 8'hA4;
                    16'h45EA: data_out = 8'hA5;
                    16'h45EB: data_out = 8'hA6;
                    16'h45EC: data_out = 8'hA7;
                    16'h45ED: data_out = 8'hA8;
                    16'h45EE: data_out = 8'hA9;
                    16'h45EF: data_out = 8'hAA;
                    16'h45F0: data_out = 8'hAB;
                    16'h45F1: data_out = 8'hAC;
                    16'h45F2: data_out = 8'hAD;
                    16'h45F3: data_out = 8'hAE;
                    16'h45F4: data_out = 8'hAF;
                    16'h45F5: data_out = 8'hB0;
                    16'h45F6: data_out = 8'hB1;
                    16'h45F7: data_out = 8'hB2;
                    16'h45F8: data_out = 8'hB3;
                    16'h45F9: data_out = 8'hB4;
                    16'h45FA: data_out = 8'hB5;
                    16'h45FB: data_out = 8'hB6;
                    16'h45FC: data_out = 8'hB7;
                    16'h45FD: data_out = 8'hB8;
                    16'h45FE: data_out = 8'hB9;
                    16'h45FF: data_out = 8'hBA;
                    16'h4600: data_out = 8'h46;
                    16'h4601: data_out = 8'h47;
                    16'h4602: data_out = 8'h48;
                    16'h4603: data_out = 8'h49;
                    16'h4604: data_out = 8'h4A;
                    16'h4605: data_out = 8'h4B;
                    16'h4606: data_out = 8'h4C;
                    16'h4607: data_out = 8'h4D;
                    16'h4608: data_out = 8'h4E;
                    16'h4609: data_out = 8'h4F;
                    16'h460A: data_out = 8'h50;
                    16'h460B: data_out = 8'h51;
                    16'h460C: data_out = 8'h52;
                    16'h460D: data_out = 8'h53;
                    16'h460E: data_out = 8'h54;
                    16'h460F: data_out = 8'h55;
                    16'h4610: data_out = 8'h56;
                    16'h4611: data_out = 8'h57;
                    16'h4612: data_out = 8'h58;
                    16'h4613: data_out = 8'h59;
                    16'h4614: data_out = 8'h5A;
                    16'h4615: data_out = 8'h5B;
                    16'h4616: data_out = 8'h5C;
                    16'h4617: data_out = 8'h5D;
                    16'h4618: data_out = 8'h5E;
                    16'h4619: data_out = 8'h5F;
                    16'h461A: data_out = 8'h60;
                    16'h461B: data_out = 8'h61;
                    16'h461C: data_out = 8'h62;
                    16'h461D: data_out = 8'h63;
                    16'h461E: data_out = 8'h64;
                    16'h461F: data_out = 8'h65;
                    16'h4620: data_out = 8'h66;
                    16'h4621: data_out = 8'h67;
                    16'h4622: data_out = 8'h68;
                    16'h4623: data_out = 8'h69;
                    16'h4624: data_out = 8'h6A;
                    16'h4625: data_out = 8'h6B;
                    16'h4626: data_out = 8'h6C;
                    16'h4627: data_out = 8'h6D;
                    16'h4628: data_out = 8'h6E;
                    16'h4629: data_out = 8'h6F;
                    16'h462A: data_out = 8'h70;
                    16'h462B: data_out = 8'h71;
                    16'h462C: data_out = 8'h72;
                    16'h462D: data_out = 8'h73;
                    16'h462E: data_out = 8'h74;
                    16'h462F: data_out = 8'h75;
                    16'h4630: data_out = 8'h76;
                    16'h4631: data_out = 8'h77;
                    16'h4632: data_out = 8'h78;
                    16'h4633: data_out = 8'h79;
                    16'h4634: data_out = 8'h7A;
                    16'h4635: data_out = 8'h7B;
                    16'h4636: data_out = 8'h7C;
                    16'h4637: data_out = 8'h7D;
                    16'h4638: data_out = 8'h7E;
                    16'h4639: data_out = 8'h7F;
                    16'h463A: data_out = 8'h80;
                    16'h463B: data_out = 8'h81;
                    16'h463C: data_out = 8'h82;
                    16'h463D: data_out = 8'h83;
                    16'h463E: data_out = 8'h84;
                    16'h463F: data_out = 8'h85;
                    16'h4640: data_out = 8'h86;
                    16'h4641: data_out = 8'h87;
                    16'h4642: data_out = 8'h88;
                    16'h4643: data_out = 8'h89;
                    16'h4644: data_out = 8'h8A;
                    16'h4645: data_out = 8'h8B;
                    16'h4646: data_out = 8'h8C;
                    16'h4647: data_out = 8'h8D;
                    16'h4648: data_out = 8'h8E;
                    16'h4649: data_out = 8'h8F;
                    16'h464A: data_out = 8'h90;
                    16'h464B: data_out = 8'h91;
                    16'h464C: data_out = 8'h92;
                    16'h464D: data_out = 8'h93;
                    16'h464E: data_out = 8'h94;
                    16'h464F: data_out = 8'h95;
                    16'h4650: data_out = 8'h96;
                    16'h4651: data_out = 8'h97;
                    16'h4652: data_out = 8'h98;
                    16'h4653: data_out = 8'h99;
                    16'h4654: data_out = 8'h9A;
                    16'h4655: data_out = 8'h9B;
                    16'h4656: data_out = 8'h9C;
                    16'h4657: data_out = 8'h9D;
                    16'h4658: data_out = 8'h9E;
                    16'h4659: data_out = 8'h9F;
                    16'h465A: data_out = 8'hA0;
                    16'h465B: data_out = 8'hA1;
                    16'h465C: data_out = 8'hA2;
                    16'h465D: data_out = 8'hA3;
                    16'h465E: data_out = 8'hA4;
                    16'h465F: data_out = 8'hA5;
                    16'h4660: data_out = 8'hA6;
                    16'h4661: data_out = 8'hA7;
                    16'h4662: data_out = 8'hA8;
                    16'h4663: data_out = 8'hA9;
                    16'h4664: data_out = 8'hAA;
                    16'h4665: data_out = 8'hAB;
                    16'h4666: data_out = 8'hAC;
                    16'h4667: data_out = 8'hAD;
                    16'h4668: data_out = 8'hAE;
                    16'h4669: data_out = 8'hAF;
                    16'h466A: data_out = 8'hB0;
                    16'h466B: data_out = 8'hB1;
                    16'h466C: data_out = 8'hB2;
                    16'h466D: data_out = 8'hB3;
                    16'h466E: data_out = 8'hB4;
                    16'h466F: data_out = 8'hB5;
                    16'h4670: data_out = 8'hB6;
                    16'h4671: data_out = 8'hB7;
                    16'h4672: data_out = 8'hB8;
                    16'h4673: data_out = 8'hB9;
                    16'h4674: data_out = 8'hBA;
                    16'h4675: data_out = 8'hBB;
                    16'h4676: data_out = 8'hBC;
                    16'h4677: data_out = 8'hBD;
                    16'h4678: data_out = 8'hBE;
                    16'h4679: data_out = 8'hBF;
                    16'h467A: data_out = 8'hC0;
                    16'h467B: data_out = 8'hC1;
                    16'h467C: data_out = 8'hC2;
                    16'h467D: data_out = 8'hC3;
                    16'h467E: data_out = 8'hC4;
                    16'h467F: data_out = 8'hC5;
                    16'h4680: data_out = 8'h46;
                    16'h4681: data_out = 8'h45;
                    16'h4682: data_out = 8'h44;
                    16'h4683: data_out = 8'h43;
                    16'h4684: data_out = 8'h42;
                    16'h4685: data_out = 8'h41;
                    16'h4686: data_out = 8'h40;
                    16'h4687: data_out = 8'h3F;
                    16'h4688: data_out = 8'h3E;
                    16'h4689: data_out = 8'h3D;
                    16'h468A: data_out = 8'h3C;
                    16'h468B: data_out = 8'h3B;
                    16'h468C: data_out = 8'h3A;
                    16'h468D: data_out = 8'h39;
                    16'h468E: data_out = 8'h38;
                    16'h468F: data_out = 8'h37;
                    16'h4690: data_out = 8'h36;
                    16'h4691: data_out = 8'h35;
                    16'h4692: data_out = 8'h34;
                    16'h4693: data_out = 8'h33;
                    16'h4694: data_out = 8'h32;
                    16'h4695: data_out = 8'h31;
                    16'h4696: data_out = 8'h30;
                    16'h4697: data_out = 8'h2F;
                    16'h4698: data_out = 8'h2E;
                    16'h4699: data_out = 8'h2D;
                    16'h469A: data_out = 8'h2C;
                    16'h469B: data_out = 8'h2B;
                    16'h469C: data_out = 8'h2A;
                    16'h469D: data_out = 8'h29;
                    16'h469E: data_out = 8'h28;
                    16'h469F: data_out = 8'h27;
                    16'h46A0: data_out = 8'h26;
                    16'h46A1: data_out = 8'h25;
                    16'h46A2: data_out = 8'h24;
                    16'h46A3: data_out = 8'h23;
                    16'h46A4: data_out = 8'h22;
                    16'h46A5: data_out = 8'h21;
                    16'h46A6: data_out = 8'h20;
                    16'h46A7: data_out = 8'h1F;
                    16'h46A8: data_out = 8'h1E;
                    16'h46A9: data_out = 8'h1D;
                    16'h46AA: data_out = 8'h1C;
                    16'h46AB: data_out = 8'h1B;
                    16'h46AC: data_out = 8'h1A;
                    16'h46AD: data_out = 8'h19;
                    16'h46AE: data_out = 8'h18;
                    16'h46AF: data_out = 8'h17;
                    16'h46B0: data_out = 8'h16;
                    16'h46B1: data_out = 8'h15;
                    16'h46B2: data_out = 8'h14;
                    16'h46B3: data_out = 8'h13;
                    16'h46B4: data_out = 8'h12;
                    16'h46B5: data_out = 8'h11;
                    16'h46B6: data_out = 8'h10;
                    16'h46B7: data_out = 8'hF;
                    16'h46B8: data_out = 8'hE;
                    16'h46B9: data_out = 8'hD;
                    16'h46BA: data_out = 8'hC;
                    16'h46BB: data_out = 8'hB;
                    16'h46BC: data_out = 8'hA;
                    16'h46BD: data_out = 8'h9;
                    16'h46BE: data_out = 8'h8;
                    16'h46BF: data_out = 8'h7;
                    16'h46C0: data_out = 8'h6;
                    16'h46C1: data_out = 8'h5;
                    16'h46C2: data_out = 8'h4;
                    16'h46C3: data_out = 8'h3;
                    16'h46C4: data_out = 8'h2;
                    16'h46C5: data_out = 8'h1;
                    16'h46C6: data_out = 8'h0;
                    16'h46C7: data_out = 8'h81;
                    16'h46C8: data_out = 8'h82;
                    16'h46C9: data_out = 8'h83;
                    16'h46CA: data_out = 8'h84;
                    16'h46CB: data_out = 8'h85;
                    16'h46CC: data_out = 8'h86;
                    16'h46CD: data_out = 8'h87;
                    16'h46CE: data_out = 8'h88;
                    16'h46CF: data_out = 8'h89;
                    16'h46D0: data_out = 8'h8A;
                    16'h46D1: data_out = 8'h8B;
                    16'h46D2: data_out = 8'h8C;
                    16'h46D3: data_out = 8'h8D;
                    16'h46D4: data_out = 8'h8E;
                    16'h46D5: data_out = 8'h8F;
                    16'h46D6: data_out = 8'h90;
                    16'h46D7: data_out = 8'h91;
                    16'h46D8: data_out = 8'h92;
                    16'h46D9: data_out = 8'h93;
                    16'h46DA: data_out = 8'h94;
                    16'h46DB: data_out = 8'h95;
                    16'h46DC: data_out = 8'h96;
                    16'h46DD: data_out = 8'h97;
                    16'h46DE: data_out = 8'h98;
                    16'h46DF: data_out = 8'h99;
                    16'h46E0: data_out = 8'h9A;
                    16'h46E1: data_out = 8'h9B;
                    16'h46E2: data_out = 8'h9C;
                    16'h46E3: data_out = 8'h9D;
                    16'h46E4: data_out = 8'h9E;
                    16'h46E5: data_out = 8'h9F;
                    16'h46E6: data_out = 8'hA0;
                    16'h46E7: data_out = 8'hA1;
                    16'h46E8: data_out = 8'hA2;
                    16'h46E9: data_out = 8'hA3;
                    16'h46EA: data_out = 8'hA4;
                    16'h46EB: data_out = 8'hA5;
                    16'h46EC: data_out = 8'hA6;
                    16'h46ED: data_out = 8'hA7;
                    16'h46EE: data_out = 8'hA8;
                    16'h46EF: data_out = 8'hA9;
                    16'h46F0: data_out = 8'hAA;
                    16'h46F1: data_out = 8'hAB;
                    16'h46F2: data_out = 8'hAC;
                    16'h46F3: data_out = 8'hAD;
                    16'h46F4: data_out = 8'hAE;
                    16'h46F5: data_out = 8'hAF;
                    16'h46F6: data_out = 8'hB0;
                    16'h46F7: data_out = 8'hB1;
                    16'h46F8: data_out = 8'hB2;
                    16'h46F9: data_out = 8'hB3;
                    16'h46FA: data_out = 8'hB4;
                    16'h46FB: data_out = 8'hB5;
                    16'h46FC: data_out = 8'hB6;
                    16'h46FD: data_out = 8'hB7;
                    16'h46FE: data_out = 8'hB8;
                    16'h46FF: data_out = 8'hB9;
                    16'h4700: data_out = 8'h47;
                    16'h4701: data_out = 8'h48;
                    16'h4702: data_out = 8'h49;
                    16'h4703: data_out = 8'h4A;
                    16'h4704: data_out = 8'h4B;
                    16'h4705: data_out = 8'h4C;
                    16'h4706: data_out = 8'h4D;
                    16'h4707: data_out = 8'h4E;
                    16'h4708: data_out = 8'h4F;
                    16'h4709: data_out = 8'h50;
                    16'h470A: data_out = 8'h51;
                    16'h470B: data_out = 8'h52;
                    16'h470C: data_out = 8'h53;
                    16'h470D: data_out = 8'h54;
                    16'h470E: data_out = 8'h55;
                    16'h470F: data_out = 8'h56;
                    16'h4710: data_out = 8'h57;
                    16'h4711: data_out = 8'h58;
                    16'h4712: data_out = 8'h59;
                    16'h4713: data_out = 8'h5A;
                    16'h4714: data_out = 8'h5B;
                    16'h4715: data_out = 8'h5C;
                    16'h4716: data_out = 8'h5D;
                    16'h4717: data_out = 8'h5E;
                    16'h4718: data_out = 8'h5F;
                    16'h4719: data_out = 8'h60;
                    16'h471A: data_out = 8'h61;
                    16'h471B: data_out = 8'h62;
                    16'h471C: data_out = 8'h63;
                    16'h471D: data_out = 8'h64;
                    16'h471E: data_out = 8'h65;
                    16'h471F: data_out = 8'h66;
                    16'h4720: data_out = 8'h67;
                    16'h4721: data_out = 8'h68;
                    16'h4722: data_out = 8'h69;
                    16'h4723: data_out = 8'h6A;
                    16'h4724: data_out = 8'h6B;
                    16'h4725: data_out = 8'h6C;
                    16'h4726: data_out = 8'h6D;
                    16'h4727: data_out = 8'h6E;
                    16'h4728: data_out = 8'h6F;
                    16'h4729: data_out = 8'h70;
                    16'h472A: data_out = 8'h71;
                    16'h472B: data_out = 8'h72;
                    16'h472C: data_out = 8'h73;
                    16'h472D: data_out = 8'h74;
                    16'h472E: data_out = 8'h75;
                    16'h472F: data_out = 8'h76;
                    16'h4730: data_out = 8'h77;
                    16'h4731: data_out = 8'h78;
                    16'h4732: data_out = 8'h79;
                    16'h4733: data_out = 8'h7A;
                    16'h4734: data_out = 8'h7B;
                    16'h4735: data_out = 8'h7C;
                    16'h4736: data_out = 8'h7D;
                    16'h4737: data_out = 8'h7E;
                    16'h4738: data_out = 8'h7F;
                    16'h4739: data_out = 8'h80;
                    16'h473A: data_out = 8'h81;
                    16'h473B: data_out = 8'h82;
                    16'h473C: data_out = 8'h83;
                    16'h473D: data_out = 8'h84;
                    16'h473E: data_out = 8'h85;
                    16'h473F: data_out = 8'h86;
                    16'h4740: data_out = 8'h87;
                    16'h4741: data_out = 8'h88;
                    16'h4742: data_out = 8'h89;
                    16'h4743: data_out = 8'h8A;
                    16'h4744: data_out = 8'h8B;
                    16'h4745: data_out = 8'h8C;
                    16'h4746: data_out = 8'h8D;
                    16'h4747: data_out = 8'h8E;
                    16'h4748: data_out = 8'h8F;
                    16'h4749: data_out = 8'h90;
                    16'h474A: data_out = 8'h91;
                    16'h474B: data_out = 8'h92;
                    16'h474C: data_out = 8'h93;
                    16'h474D: data_out = 8'h94;
                    16'h474E: data_out = 8'h95;
                    16'h474F: data_out = 8'h96;
                    16'h4750: data_out = 8'h97;
                    16'h4751: data_out = 8'h98;
                    16'h4752: data_out = 8'h99;
                    16'h4753: data_out = 8'h9A;
                    16'h4754: data_out = 8'h9B;
                    16'h4755: data_out = 8'h9C;
                    16'h4756: data_out = 8'h9D;
                    16'h4757: data_out = 8'h9E;
                    16'h4758: data_out = 8'h9F;
                    16'h4759: data_out = 8'hA0;
                    16'h475A: data_out = 8'hA1;
                    16'h475B: data_out = 8'hA2;
                    16'h475C: data_out = 8'hA3;
                    16'h475D: data_out = 8'hA4;
                    16'h475E: data_out = 8'hA5;
                    16'h475F: data_out = 8'hA6;
                    16'h4760: data_out = 8'hA7;
                    16'h4761: data_out = 8'hA8;
                    16'h4762: data_out = 8'hA9;
                    16'h4763: data_out = 8'hAA;
                    16'h4764: data_out = 8'hAB;
                    16'h4765: data_out = 8'hAC;
                    16'h4766: data_out = 8'hAD;
                    16'h4767: data_out = 8'hAE;
                    16'h4768: data_out = 8'hAF;
                    16'h4769: data_out = 8'hB0;
                    16'h476A: data_out = 8'hB1;
                    16'h476B: data_out = 8'hB2;
                    16'h476C: data_out = 8'hB3;
                    16'h476D: data_out = 8'hB4;
                    16'h476E: data_out = 8'hB5;
                    16'h476F: data_out = 8'hB6;
                    16'h4770: data_out = 8'hB7;
                    16'h4771: data_out = 8'hB8;
                    16'h4772: data_out = 8'hB9;
                    16'h4773: data_out = 8'hBA;
                    16'h4774: data_out = 8'hBB;
                    16'h4775: data_out = 8'hBC;
                    16'h4776: data_out = 8'hBD;
                    16'h4777: data_out = 8'hBE;
                    16'h4778: data_out = 8'hBF;
                    16'h4779: data_out = 8'hC0;
                    16'h477A: data_out = 8'hC1;
                    16'h477B: data_out = 8'hC2;
                    16'h477C: data_out = 8'hC3;
                    16'h477D: data_out = 8'hC4;
                    16'h477E: data_out = 8'hC5;
                    16'h477F: data_out = 8'hC6;
                    16'h4780: data_out = 8'h47;
                    16'h4781: data_out = 8'h46;
                    16'h4782: data_out = 8'h45;
                    16'h4783: data_out = 8'h44;
                    16'h4784: data_out = 8'h43;
                    16'h4785: data_out = 8'h42;
                    16'h4786: data_out = 8'h41;
                    16'h4787: data_out = 8'h40;
                    16'h4788: data_out = 8'h3F;
                    16'h4789: data_out = 8'h3E;
                    16'h478A: data_out = 8'h3D;
                    16'h478B: data_out = 8'h3C;
                    16'h478C: data_out = 8'h3B;
                    16'h478D: data_out = 8'h3A;
                    16'h478E: data_out = 8'h39;
                    16'h478F: data_out = 8'h38;
                    16'h4790: data_out = 8'h37;
                    16'h4791: data_out = 8'h36;
                    16'h4792: data_out = 8'h35;
                    16'h4793: data_out = 8'h34;
                    16'h4794: data_out = 8'h33;
                    16'h4795: data_out = 8'h32;
                    16'h4796: data_out = 8'h31;
                    16'h4797: data_out = 8'h30;
                    16'h4798: data_out = 8'h2F;
                    16'h4799: data_out = 8'h2E;
                    16'h479A: data_out = 8'h2D;
                    16'h479B: data_out = 8'h2C;
                    16'h479C: data_out = 8'h2B;
                    16'h479D: data_out = 8'h2A;
                    16'h479E: data_out = 8'h29;
                    16'h479F: data_out = 8'h28;
                    16'h47A0: data_out = 8'h27;
                    16'h47A1: data_out = 8'h26;
                    16'h47A2: data_out = 8'h25;
                    16'h47A3: data_out = 8'h24;
                    16'h47A4: data_out = 8'h23;
                    16'h47A5: data_out = 8'h22;
                    16'h47A6: data_out = 8'h21;
                    16'h47A7: data_out = 8'h20;
                    16'h47A8: data_out = 8'h1F;
                    16'h47A9: data_out = 8'h1E;
                    16'h47AA: data_out = 8'h1D;
                    16'h47AB: data_out = 8'h1C;
                    16'h47AC: data_out = 8'h1B;
                    16'h47AD: data_out = 8'h1A;
                    16'h47AE: data_out = 8'h19;
                    16'h47AF: data_out = 8'h18;
                    16'h47B0: data_out = 8'h17;
                    16'h47B1: data_out = 8'h16;
                    16'h47B2: data_out = 8'h15;
                    16'h47B3: data_out = 8'h14;
                    16'h47B4: data_out = 8'h13;
                    16'h47B5: data_out = 8'h12;
                    16'h47B6: data_out = 8'h11;
                    16'h47B7: data_out = 8'h10;
                    16'h47B8: data_out = 8'hF;
                    16'h47B9: data_out = 8'hE;
                    16'h47BA: data_out = 8'hD;
                    16'h47BB: data_out = 8'hC;
                    16'h47BC: data_out = 8'hB;
                    16'h47BD: data_out = 8'hA;
                    16'h47BE: data_out = 8'h9;
                    16'h47BF: data_out = 8'h8;
                    16'h47C0: data_out = 8'h7;
                    16'h47C1: data_out = 8'h6;
                    16'h47C2: data_out = 8'h5;
                    16'h47C3: data_out = 8'h4;
                    16'h47C4: data_out = 8'h3;
                    16'h47C5: data_out = 8'h2;
                    16'h47C6: data_out = 8'h1;
                    16'h47C7: data_out = 8'h0;
                    16'h47C8: data_out = 8'h81;
                    16'h47C9: data_out = 8'h82;
                    16'h47CA: data_out = 8'h83;
                    16'h47CB: data_out = 8'h84;
                    16'h47CC: data_out = 8'h85;
                    16'h47CD: data_out = 8'h86;
                    16'h47CE: data_out = 8'h87;
                    16'h47CF: data_out = 8'h88;
                    16'h47D0: data_out = 8'h89;
                    16'h47D1: data_out = 8'h8A;
                    16'h47D2: data_out = 8'h8B;
                    16'h47D3: data_out = 8'h8C;
                    16'h47D4: data_out = 8'h8D;
                    16'h47D5: data_out = 8'h8E;
                    16'h47D6: data_out = 8'h8F;
                    16'h47D7: data_out = 8'h90;
                    16'h47D8: data_out = 8'h91;
                    16'h47D9: data_out = 8'h92;
                    16'h47DA: data_out = 8'h93;
                    16'h47DB: data_out = 8'h94;
                    16'h47DC: data_out = 8'h95;
                    16'h47DD: data_out = 8'h96;
                    16'h47DE: data_out = 8'h97;
                    16'h47DF: data_out = 8'h98;
                    16'h47E0: data_out = 8'h99;
                    16'h47E1: data_out = 8'h9A;
                    16'h47E2: data_out = 8'h9B;
                    16'h47E3: data_out = 8'h9C;
                    16'h47E4: data_out = 8'h9D;
                    16'h47E5: data_out = 8'h9E;
                    16'h47E6: data_out = 8'h9F;
                    16'h47E7: data_out = 8'hA0;
                    16'h47E8: data_out = 8'hA1;
                    16'h47E9: data_out = 8'hA2;
                    16'h47EA: data_out = 8'hA3;
                    16'h47EB: data_out = 8'hA4;
                    16'h47EC: data_out = 8'hA5;
                    16'h47ED: data_out = 8'hA6;
                    16'h47EE: data_out = 8'hA7;
                    16'h47EF: data_out = 8'hA8;
                    16'h47F0: data_out = 8'hA9;
                    16'h47F1: data_out = 8'hAA;
                    16'h47F2: data_out = 8'hAB;
                    16'h47F3: data_out = 8'hAC;
                    16'h47F4: data_out = 8'hAD;
                    16'h47F5: data_out = 8'hAE;
                    16'h47F6: data_out = 8'hAF;
                    16'h47F7: data_out = 8'hB0;
                    16'h47F8: data_out = 8'hB1;
                    16'h47F9: data_out = 8'hB2;
                    16'h47FA: data_out = 8'hB3;
                    16'h47FB: data_out = 8'hB4;
                    16'h47FC: data_out = 8'hB5;
                    16'h47FD: data_out = 8'hB6;
                    16'h47FE: data_out = 8'hB7;
                    16'h47FF: data_out = 8'hB8;
                    16'h4800: data_out = 8'h48;
                    16'h4801: data_out = 8'h49;
                    16'h4802: data_out = 8'h4A;
                    16'h4803: data_out = 8'h4B;
                    16'h4804: data_out = 8'h4C;
                    16'h4805: data_out = 8'h4D;
                    16'h4806: data_out = 8'h4E;
                    16'h4807: data_out = 8'h4F;
                    16'h4808: data_out = 8'h50;
                    16'h4809: data_out = 8'h51;
                    16'h480A: data_out = 8'h52;
                    16'h480B: data_out = 8'h53;
                    16'h480C: data_out = 8'h54;
                    16'h480D: data_out = 8'h55;
                    16'h480E: data_out = 8'h56;
                    16'h480F: data_out = 8'h57;
                    16'h4810: data_out = 8'h58;
                    16'h4811: data_out = 8'h59;
                    16'h4812: data_out = 8'h5A;
                    16'h4813: data_out = 8'h5B;
                    16'h4814: data_out = 8'h5C;
                    16'h4815: data_out = 8'h5D;
                    16'h4816: data_out = 8'h5E;
                    16'h4817: data_out = 8'h5F;
                    16'h4818: data_out = 8'h60;
                    16'h4819: data_out = 8'h61;
                    16'h481A: data_out = 8'h62;
                    16'h481B: data_out = 8'h63;
                    16'h481C: data_out = 8'h64;
                    16'h481D: data_out = 8'h65;
                    16'h481E: data_out = 8'h66;
                    16'h481F: data_out = 8'h67;
                    16'h4820: data_out = 8'h68;
                    16'h4821: data_out = 8'h69;
                    16'h4822: data_out = 8'h6A;
                    16'h4823: data_out = 8'h6B;
                    16'h4824: data_out = 8'h6C;
                    16'h4825: data_out = 8'h6D;
                    16'h4826: data_out = 8'h6E;
                    16'h4827: data_out = 8'h6F;
                    16'h4828: data_out = 8'h70;
                    16'h4829: data_out = 8'h71;
                    16'h482A: data_out = 8'h72;
                    16'h482B: data_out = 8'h73;
                    16'h482C: data_out = 8'h74;
                    16'h482D: data_out = 8'h75;
                    16'h482E: data_out = 8'h76;
                    16'h482F: data_out = 8'h77;
                    16'h4830: data_out = 8'h78;
                    16'h4831: data_out = 8'h79;
                    16'h4832: data_out = 8'h7A;
                    16'h4833: data_out = 8'h7B;
                    16'h4834: data_out = 8'h7C;
                    16'h4835: data_out = 8'h7D;
                    16'h4836: data_out = 8'h7E;
                    16'h4837: data_out = 8'h7F;
                    16'h4838: data_out = 8'h80;
                    16'h4839: data_out = 8'h81;
                    16'h483A: data_out = 8'h82;
                    16'h483B: data_out = 8'h83;
                    16'h483C: data_out = 8'h84;
                    16'h483D: data_out = 8'h85;
                    16'h483E: data_out = 8'h86;
                    16'h483F: data_out = 8'h87;
                    16'h4840: data_out = 8'h88;
                    16'h4841: data_out = 8'h89;
                    16'h4842: data_out = 8'h8A;
                    16'h4843: data_out = 8'h8B;
                    16'h4844: data_out = 8'h8C;
                    16'h4845: data_out = 8'h8D;
                    16'h4846: data_out = 8'h8E;
                    16'h4847: data_out = 8'h8F;
                    16'h4848: data_out = 8'h90;
                    16'h4849: data_out = 8'h91;
                    16'h484A: data_out = 8'h92;
                    16'h484B: data_out = 8'h93;
                    16'h484C: data_out = 8'h94;
                    16'h484D: data_out = 8'h95;
                    16'h484E: data_out = 8'h96;
                    16'h484F: data_out = 8'h97;
                    16'h4850: data_out = 8'h98;
                    16'h4851: data_out = 8'h99;
                    16'h4852: data_out = 8'h9A;
                    16'h4853: data_out = 8'h9B;
                    16'h4854: data_out = 8'h9C;
                    16'h4855: data_out = 8'h9D;
                    16'h4856: data_out = 8'h9E;
                    16'h4857: data_out = 8'h9F;
                    16'h4858: data_out = 8'hA0;
                    16'h4859: data_out = 8'hA1;
                    16'h485A: data_out = 8'hA2;
                    16'h485B: data_out = 8'hA3;
                    16'h485C: data_out = 8'hA4;
                    16'h485D: data_out = 8'hA5;
                    16'h485E: data_out = 8'hA6;
                    16'h485F: data_out = 8'hA7;
                    16'h4860: data_out = 8'hA8;
                    16'h4861: data_out = 8'hA9;
                    16'h4862: data_out = 8'hAA;
                    16'h4863: data_out = 8'hAB;
                    16'h4864: data_out = 8'hAC;
                    16'h4865: data_out = 8'hAD;
                    16'h4866: data_out = 8'hAE;
                    16'h4867: data_out = 8'hAF;
                    16'h4868: data_out = 8'hB0;
                    16'h4869: data_out = 8'hB1;
                    16'h486A: data_out = 8'hB2;
                    16'h486B: data_out = 8'hB3;
                    16'h486C: data_out = 8'hB4;
                    16'h486D: data_out = 8'hB5;
                    16'h486E: data_out = 8'hB6;
                    16'h486F: data_out = 8'hB7;
                    16'h4870: data_out = 8'hB8;
                    16'h4871: data_out = 8'hB9;
                    16'h4872: data_out = 8'hBA;
                    16'h4873: data_out = 8'hBB;
                    16'h4874: data_out = 8'hBC;
                    16'h4875: data_out = 8'hBD;
                    16'h4876: data_out = 8'hBE;
                    16'h4877: data_out = 8'hBF;
                    16'h4878: data_out = 8'hC0;
                    16'h4879: data_out = 8'hC1;
                    16'h487A: data_out = 8'hC2;
                    16'h487B: data_out = 8'hC3;
                    16'h487C: data_out = 8'hC4;
                    16'h487D: data_out = 8'hC5;
                    16'h487E: data_out = 8'hC6;
                    16'h487F: data_out = 8'hC7;
                    16'h4880: data_out = 8'h48;
                    16'h4881: data_out = 8'h47;
                    16'h4882: data_out = 8'h46;
                    16'h4883: data_out = 8'h45;
                    16'h4884: data_out = 8'h44;
                    16'h4885: data_out = 8'h43;
                    16'h4886: data_out = 8'h42;
                    16'h4887: data_out = 8'h41;
                    16'h4888: data_out = 8'h40;
                    16'h4889: data_out = 8'h3F;
                    16'h488A: data_out = 8'h3E;
                    16'h488B: data_out = 8'h3D;
                    16'h488C: data_out = 8'h3C;
                    16'h488D: data_out = 8'h3B;
                    16'h488E: data_out = 8'h3A;
                    16'h488F: data_out = 8'h39;
                    16'h4890: data_out = 8'h38;
                    16'h4891: data_out = 8'h37;
                    16'h4892: data_out = 8'h36;
                    16'h4893: data_out = 8'h35;
                    16'h4894: data_out = 8'h34;
                    16'h4895: data_out = 8'h33;
                    16'h4896: data_out = 8'h32;
                    16'h4897: data_out = 8'h31;
                    16'h4898: data_out = 8'h30;
                    16'h4899: data_out = 8'h2F;
                    16'h489A: data_out = 8'h2E;
                    16'h489B: data_out = 8'h2D;
                    16'h489C: data_out = 8'h2C;
                    16'h489D: data_out = 8'h2B;
                    16'h489E: data_out = 8'h2A;
                    16'h489F: data_out = 8'h29;
                    16'h48A0: data_out = 8'h28;
                    16'h48A1: data_out = 8'h27;
                    16'h48A2: data_out = 8'h26;
                    16'h48A3: data_out = 8'h25;
                    16'h48A4: data_out = 8'h24;
                    16'h48A5: data_out = 8'h23;
                    16'h48A6: data_out = 8'h22;
                    16'h48A7: data_out = 8'h21;
                    16'h48A8: data_out = 8'h20;
                    16'h48A9: data_out = 8'h1F;
                    16'h48AA: data_out = 8'h1E;
                    16'h48AB: data_out = 8'h1D;
                    16'h48AC: data_out = 8'h1C;
                    16'h48AD: data_out = 8'h1B;
                    16'h48AE: data_out = 8'h1A;
                    16'h48AF: data_out = 8'h19;
                    16'h48B0: data_out = 8'h18;
                    16'h48B1: data_out = 8'h17;
                    16'h48B2: data_out = 8'h16;
                    16'h48B3: data_out = 8'h15;
                    16'h48B4: data_out = 8'h14;
                    16'h48B5: data_out = 8'h13;
                    16'h48B6: data_out = 8'h12;
                    16'h48B7: data_out = 8'h11;
                    16'h48B8: data_out = 8'h10;
                    16'h48B9: data_out = 8'hF;
                    16'h48BA: data_out = 8'hE;
                    16'h48BB: data_out = 8'hD;
                    16'h48BC: data_out = 8'hC;
                    16'h48BD: data_out = 8'hB;
                    16'h48BE: data_out = 8'hA;
                    16'h48BF: data_out = 8'h9;
                    16'h48C0: data_out = 8'h8;
                    16'h48C1: data_out = 8'h7;
                    16'h48C2: data_out = 8'h6;
                    16'h48C3: data_out = 8'h5;
                    16'h48C4: data_out = 8'h4;
                    16'h48C5: data_out = 8'h3;
                    16'h48C6: data_out = 8'h2;
                    16'h48C7: data_out = 8'h1;
                    16'h48C8: data_out = 8'h0;
                    16'h48C9: data_out = 8'h81;
                    16'h48CA: data_out = 8'h82;
                    16'h48CB: data_out = 8'h83;
                    16'h48CC: data_out = 8'h84;
                    16'h48CD: data_out = 8'h85;
                    16'h48CE: data_out = 8'h86;
                    16'h48CF: data_out = 8'h87;
                    16'h48D0: data_out = 8'h88;
                    16'h48D1: data_out = 8'h89;
                    16'h48D2: data_out = 8'h8A;
                    16'h48D3: data_out = 8'h8B;
                    16'h48D4: data_out = 8'h8C;
                    16'h48D5: data_out = 8'h8D;
                    16'h48D6: data_out = 8'h8E;
                    16'h48D7: data_out = 8'h8F;
                    16'h48D8: data_out = 8'h90;
                    16'h48D9: data_out = 8'h91;
                    16'h48DA: data_out = 8'h92;
                    16'h48DB: data_out = 8'h93;
                    16'h48DC: data_out = 8'h94;
                    16'h48DD: data_out = 8'h95;
                    16'h48DE: data_out = 8'h96;
                    16'h48DF: data_out = 8'h97;
                    16'h48E0: data_out = 8'h98;
                    16'h48E1: data_out = 8'h99;
                    16'h48E2: data_out = 8'h9A;
                    16'h48E3: data_out = 8'h9B;
                    16'h48E4: data_out = 8'h9C;
                    16'h48E5: data_out = 8'h9D;
                    16'h48E6: data_out = 8'h9E;
                    16'h48E7: data_out = 8'h9F;
                    16'h48E8: data_out = 8'hA0;
                    16'h48E9: data_out = 8'hA1;
                    16'h48EA: data_out = 8'hA2;
                    16'h48EB: data_out = 8'hA3;
                    16'h48EC: data_out = 8'hA4;
                    16'h48ED: data_out = 8'hA5;
                    16'h48EE: data_out = 8'hA6;
                    16'h48EF: data_out = 8'hA7;
                    16'h48F0: data_out = 8'hA8;
                    16'h48F1: data_out = 8'hA9;
                    16'h48F2: data_out = 8'hAA;
                    16'h48F3: data_out = 8'hAB;
                    16'h48F4: data_out = 8'hAC;
                    16'h48F5: data_out = 8'hAD;
                    16'h48F6: data_out = 8'hAE;
                    16'h48F7: data_out = 8'hAF;
                    16'h48F8: data_out = 8'hB0;
                    16'h48F9: data_out = 8'hB1;
                    16'h48FA: data_out = 8'hB2;
                    16'h48FB: data_out = 8'hB3;
                    16'h48FC: data_out = 8'hB4;
                    16'h48FD: data_out = 8'hB5;
                    16'h48FE: data_out = 8'hB6;
                    16'h48FF: data_out = 8'hB7;
                    16'h4900: data_out = 8'h49;
                    16'h4901: data_out = 8'h4A;
                    16'h4902: data_out = 8'h4B;
                    16'h4903: data_out = 8'h4C;
                    16'h4904: data_out = 8'h4D;
                    16'h4905: data_out = 8'h4E;
                    16'h4906: data_out = 8'h4F;
                    16'h4907: data_out = 8'h50;
                    16'h4908: data_out = 8'h51;
                    16'h4909: data_out = 8'h52;
                    16'h490A: data_out = 8'h53;
                    16'h490B: data_out = 8'h54;
                    16'h490C: data_out = 8'h55;
                    16'h490D: data_out = 8'h56;
                    16'h490E: data_out = 8'h57;
                    16'h490F: data_out = 8'h58;
                    16'h4910: data_out = 8'h59;
                    16'h4911: data_out = 8'h5A;
                    16'h4912: data_out = 8'h5B;
                    16'h4913: data_out = 8'h5C;
                    16'h4914: data_out = 8'h5D;
                    16'h4915: data_out = 8'h5E;
                    16'h4916: data_out = 8'h5F;
                    16'h4917: data_out = 8'h60;
                    16'h4918: data_out = 8'h61;
                    16'h4919: data_out = 8'h62;
                    16'h491A: data_out = 8'h63;
                    16'h491B: data_out = 8'h64;
                    16'h491C: data_out = 8'h65;
                    16'h491D: data_out = 8'h66;
                    16'h491E: data_out = 8'h67;
                    16'h491F: data_out = 8'h68;
                    16'h4920: data_out = 8'h69;
                    16'h4921: data_out = 8'h6A;
                    16'h4922: data_out = 8'h6B;
                    16'h4923: data_out = 8'h6C;
                    16'h4924: data_out = 8'h6D;
                    16'h4925: data_out = 8'h6E;
                    16'h4926: data_out = 8'h6F;
                    16'h4927: data_out = 8'h70;
                    16'h4928: data_out = 8'h71;
                    16'h4929: data_out = 8'h72;
                    16'h492A: data_out = 8'h73;
                    16'h492B: data_out = 8'h74;
                    16'h492C: data_out = 8'h75;
                    16'h492D: data_out = 8'h76;
                    16'h492E: data_out = 8'h77;
                    16'h492F: data_out = 8'h78;
                    16'h4930: data_out = 8'h79;
                    16'h4931: data_out = 8'h7A;
                    16'h4932: data_out = 8'h7B;
                    16'h4933: data_out = 8'h7C;
                    16'h4934: data_out = 8'h7D;
                    16'h4935: data_out = 8'h7E;
                    16'h4936: data_out = 8'h7F;
                    16'h4937: data_out = 8'h80;
                    16'h4938: data_out = 8'h81;
                    16'h4939: data_out = 8'h82;
                    16'h493A: data_out = 8'h83;
                    16'h493B: data_out = 8'h84;
                    16'h493C: data_out = 8'h85;
                    16'h493D: data_out = 8'h86;
                    16'h493E: data_out = 8'h87;
                    16'h493F: data_out = 8'h88;
                    16'h4940: data_out = 8'h89;
                    16'h4941: data_out = 8'h8A;
                    16'h4942: data_out = 8'h8B;
                    16'h4943: data_out = 8'h8C;
                    16'h4944: data_out = 8'h8D;
                    16'h4945: data_out = 8'h8E;
                    16'h4946: data_out = 8'h8F;
                    16'h4947: data_out = 8'h90;
                    16'h4948: data_out = 8'h91;
                    16'h4949: data_out = 8'h92;
                    16'h494A: data_out = 8'h93;
                    16'h494B: data_out = 8'h94;
                    16'h494C: data_out = 8'h95;
                    16'h494D: data_out = 8'h96;
                    16'h494E: data_out = 8'h97;
                    16'h494F: data_out = 8'h98;
                    16'h4950: data_out = 8'h99;
                    16'h4951: data_out = 8'h9A;
                    16'h4952: data_out = 8'h9B;
                    16'h4953: data_out = 8'h9C;
                    16'h4954: data_out = 8'h9D;
                    16'h4955: data_out = 8'h9E;
                    16'h4956: data_out = 8'h9F;
                    16'h4957: data_out = 8'hA0;
                    16'h4958: data_out = 8'hA1;
                    16'h4959: data_out = 8'hA2;
                    16'h495A: data_out = 8'hA3;
                    16'h495B: data_out = 8'hA4;
                    16'h495C: data_out = 8'hA5;
                    16'h495D: data_out = 8'hA6;
                    16'h495E: data_out = 8'hA7;
                    16'h495F: data_out = 8'hA8;
                    16'h4960: data_out = 8'hA9;
                    16'h4961: data_out = 8'hAA;
                    16'h4962: data_out = 8'hAB;
                    16'h4963: data_out = 8'hAC;
                    16'h4964: data_out = 8'hAD;
                    16'h4965: data_out = 8'hAE;
                    16'h4966: data_out = 8'hAF;
                    16'h4967: data_out = 8'hB0;
                    16'h4968: data_out = 8'hB1;
                    16'h4969: data_out = 8'hB2;
                    16'h496A: data_out = 8'hB3;
                    16'h496B: data_out = 8'hB4;
                    16'h496C: data_out = 8'hB5;
                    16'h496D: data_out = 8'hB6;
                    16'h496E: data_out = 8'hB7;
                    16'h496F: data_out = 8'hB8;
                    16'h4970: data_out = 8'hB9;
                    16'h4971: data_out = 8'hBA;
                    16'h4972: data_out = 8'hBB;
                    16'h4973: data_out = 8'hBC;
                    16'h4974: data_out = 8'hBD;
                    16'h4975: data_out = 8'hBE;
                    16'h4976: data_out = 8'hBF;
                    16'h4977: data_out = 8'hC0;
                    16'h4978: data_out = 8'hC1;
                    16'h4979: data_out = 8'hC2;
                    16'h497A: data_out = 8'hC3;
                    16'h497B: data_out = 8'hC4;
                    16'h497C: data_out = 8'hC5;
                    16'h497D: data_out = 8'hC6;
                    16'h497E: data_out = 8'hC7;
                    16'h497F: data_out = 8'hC8;
                    16'h4980: data_out = 8'h49;
                    16'h4981: data_out = 8'h48;
                    16'h4982: data_out = 8'h47;
                    16'h4983: data_out = 8'h46;
                    16'h4984: data_out = 8'h45;
                    16'h4985: data_out = 8'h44;
                    16'h4986: data_out = 8'h43;
                    16'h4987: data_out = 8'h42;
                    16'h4988: data_out = 8'h41;
                    16'h4989: data_out = 8'h40;
                    16'h498A: data_out = 8'h3F;
                    16'h498B: data_out = 8'h3E;
                    16'h498C: data_out = 8'h3D;
                    16'h498D: data_out = 8'h3C;
                    16'h498E: data_out = 8'h3B;
                    16'h498F: data_out = 8'h3A;
                    16'h4990: data_out = 8'h39;
                    16'h4991: data_out = 8'h38;
                    16'h4992: data_out = 8'h37;
                    16'h4993: data_out = 8'h36;
                    16'h4994: data_out = 8'h35;
                    16'h4995: data_out = 8'h34;
                    16'h4996: data_out = 8'h33;
                    16'h4997: data_out = 8'h32;
                    16'h4998: data_out = 8'h31;
                    16'h4999: data_out = 8'h30;
                    16'h499A: data_out = 8'h2F;
                    16'h499B: data_out = 8'h2E;
                    16'h499C: data_out = 8'h2D;
                    16'h499D: data_out = 8'h2C;
                    16'h499E: data_out = 8'h2B;
                    16'h499F: data_out = 8'h2A;
                    16'h49A0: data_out = 8'h29;
                    16'h49A1: data_out = 8'h28;
                    16'h49A2: data_out = 8'h27;
                    16'h49A3: data_out = 8'h26;
                    16'h49A4: data_out = 8'h25;
                    16'h49A5: data_out = 8'h24;
                    16'h49A6: data_out = 8'h23;
                    16'h49A7: data_out = 8'h22;
                    16'h49A8: data_out = 8'h21;
                    16'h49A9: data_out = 8'h20;
                    16'h49AA: data_out = 8'h1F;
                    16'h49AB: data_out = 8'h1E;
                    16'h49AC: data_out = 8'h1D;
                    16'h49AD: data_out = 8'h1C;
                    16'h49AE: data_out = 8'h1B;
                    16'h49AF: data_out = 8'h1A;
                    16'h49B0: data_out = 8'h19;
                    16'h49B1: data_out = 8'h18;
                    16'h49B2: data_out = 8'h17;
                    16'h49B3: data_out = 8'h16;
                    16'h49B4: data_out = 8'h15;
                    16'h49B5: data_out = 8'h14;
                    16'h49B6: data_out = 8'h13;
                    16'h49B7: data_out = 8'h12;
                    16'h49B8: data_out = 8'h11;
                    16'h49B9: data_out = 8'h10;
                    16'h49BA: data_out = 8'hF;
                    16'h49BB: data_out = 8'hE;
                    16'h49BC: data_out = 8'hD;
                    16'h49BD: data_out = 8'hC;
                    16'h49BE: data_out = 8'hB;
                    16'h49BF: data_out = 8'hA;
                    16'h49C0: data_out = 8'h9;
                    16'h49C1: data_out = 8'h8;
                    16'h49C2: data_out = 8'h7;
                    16'h49C3: data_out = 8'h6;
                    16'h49C4: data_out = 8'h5;
                    16'h49C5: data_out = 8'h4;
                    16'h49C6: data_out = 8'h3;
                    16'h49C7: data_out = 8'h2;
                    16'h49C8: data_out = 8'h1;
                    16'h49C9: data_out = 8'h0;
                    16'h49CA: data_out = 8'h81;
                    16'h49CB: data_out = 8'h82;
                    16'h49CC: data_out = 8'h83;
                    16'h49CD: data_out = 8'h84;
                    16'h49CE: data_out = 8'h85;
                    16'h49CF: data_out = 8'h86;
                    16'h49D0: data_out = 8'h87;
                    16'h49D1: data_out = 8'h88;
                    16'h49D2: data_out = 8'h89;
                    16'h49D3: data_out = 8'h8A;
                    16'h49D4: data_out = 8'h8B;
                    16'h49D5: data_out = 8'h8C;
                    16'h49D6: data_out = 8'h8D;
                    16'h49D7: data_out = 8'h8E;
                    16'h49D8: data_out = 8'h8F;
                    16'h49D9: data_out = 8'h90;
                    16'h49DA: data_out = 8'h91;
                    16'h49DB: data_out = 8'h92;
                    16'h49DC: data_out = 8'h93;
                    16'h49DD: data_out = 8'h94;
                    16'h49DE: data_out = 8'h95;
                    16'h49DF: data_out = 8'h96;
                    16'h49E0: data_out = 8'h97;
                    16'h49E1: data_out = 8'h98;
                    16'h49E2: data_out = 8'h99;
                    16'h49E3: data_out = 8'h9A;
                    16'h49E4: data_out = 8'h9B;
                    16'h49E5: data_out = 8'h9C;
                    16'h49E6: data_out = 8'h9D;
                    16'h49E7: data_out = 8'h9E;
                    16'h49E8: data_out = 8'h9F;
                    16'h49E9: data_out = 8'hA0;
                    16'h49EA: data_out = 8'hA1;
                    16'h49EB: data_out = 8'hA2;
                    16'h49EC: data_out = 8'hA3;
                    16'h49ED: data_out = 8'hA4;
                    16'h49EE: data_out = 8'hA5;
                    16'h49EF: data_out = 8'hA6;
                    16'h49F0: data_out = 8'hA7;
                    16'h49F1: data_out = 8'hA8;
                    16'h49F2: data_out = 8'hA9;
                    16'h49F3: data_out = 8'hAA;
                    16'h49F4: data_out = 8'hAB;
                    16'h49F5: data_out = 8'hAC;
                    16'h49F6: data_out = 8'hAD;
                    16'h49F7: data_out = 8'hAE;
                    16'h49F8: data_out = 8'hAF;
                    16'h49F9: data_out = 8'hB0;
                    16'h49FA: data_out = 8'hB1;
                    16'h49FB: data_out = 8'hB2;
                    16'h49FC: data_out = 8'hB3;
                    16'h49FD: data_out = 8'hB4;
                    16'h49FE: data_out = 8'hB5;
                    16'h49FF: data_out = 8'hB6;
                    16'h4A00: data_out = 8'h4A;
                    16'h4A01: data_out = 8'h4B;
                    16'h4A02: data_out = 8'h4C;
                    16'h4A03: data_out = 8'h4D;
                    16'h4A04: data_out = 8'h4E;
                    16'h4A05: data_out = 8'h4F;
                    16'h4A06: data_out = 8'h50;
                    16'h4A07: data_out = 8'h51;
                    16'h4A08: data_out = 8'h52;
                    16'h4A09: data_out = 8'h53;
                    16'h4A0A: data_out = 8'h54;
                    16'h4A0B: data_out = 8'h55;
                    16'h4A0C: data_out = 8'h56;
                    16'h4A0D: data_out = 8'h57;
                    16'h4A0E: data_out = 8'h58;
                    16'h4A0F: data_out = 8'h59;
                    16'h4A10: data_out = 8'h5A;
                    16'h4A11: data_out = 8'h5B;
                    16'h4A12: data_out = 8'h5C;
                    16'h4A13: data_out = 8'h5D;
                    16'h4A14: data_out = 8'h5E;
                    16'h4A15: data_out = 8'h5F;
                    16'h4A16: data_out = 8'h60;
                    16'h4A17: data_out = 8'h61;
                    16'h4A18: data_out = 8'h62;
                    16'h4A19: data_out = 8'h63;
                    16'h4A1A: data_out = 8'h64;
                    16'h4A1B: data_out = 8'h65;
                    16'h4A1C: data_out = 8'h66;
                    16'h4A1D: data_out = 8'h67;
                    16'h4A1E: data_out = 8'h68;
                    16'h4A1F: data_out = 8'h69;
                    16'h4A20: data_out = 8'h6A;
                    16'h4A21: data_out = 8'h6B;
                    16'h4A22: data_out = 8'h6C;
                    16'h4A23: data_out = 8'h6D;
                    16'h4A24: data_out = 8'h6E;
                    16'h4A25: data_out = 8'h6F;
                    16'h4A26: data_out = 8'h70;
                    16'h4A27: data_out = 8'h71;
                    16'h4A28: data_out = 8'h72;
                    16'h4A29: data_out = 8'h73;
                    16'h4A2A: data_out = 8'h74;
                    16'h4A2B: data_out = 8'h75;
                    16'h4A2C: data_out = 8'h76;
                    16'h4A2D: data_out = 8'h77;
                    16'h4A2E: data_out = 8'h78;
                    16'h4A2F: data_out = 8'h79;
                    16'h4A30: data_out = 8'h7A;
                    16'h4A31: data_out = 8'h7B;
                    16'h4A32: data_out = 8'h7C;
                    16'h4A33: data_out = 8'h7D;
                    16'h4A34: data_out = 8'h7E;
                    16'h4A35: data_out = 8'h7F;
                    16'h4A36: data_out = 8'h80;
                    16'h4A37: data_out = 8'h81;
                    16'h4A38: data_out = 8'h82;
                    16'h4A39: data_out = 8'h83;
                    16'h4A3A: data_out = 8'h84;
                    16'h4A3B: data_out = 8'h85;
                    16'h4A3C: data_out = 8'h86;
                    16'h4A3D: data_out = 8'h87;
                    16'h4A3E: data_out = 8'h88;
                    16'h4A3F: data_out = 8'h89;
                    16'h4A40: data_out = 8'h8A;
                    16'h4A41: data_out = 8'h8B;
                    16'h4A42: data_out = 8'h8C;
                    16'h4A43: data_out = 8'h8D;
                    16'h4A44: data_out = 8'h8E;
                    16'h4A45: data_out = 8'h8F;
                    16'h4A46: data_out = 8'h90;
                    16'h4A47: data_out = 8'h91;
                    16'h4A48: data_out = 8'h92;
                    16'h4A49: data_out = 8'h93;
                    16'h4A4A: data_out = 8'h94;
                    16'h4A4B: data_out = 8'h95;
                    16'h4A4C: data_out = 8'h96;
                    16'h4A4D: data_out = 8'h97;
                    16'h4A4E: data_out = 8'h98;
                    16'h4A4F: data_out = 8'h99;
                    16'h4A50: data_out = 8'h9A;
                    16'h4A51: data_out = 8'h9B;
                    16'h4A52: data_out = 8'h9C;
                    16'h4A53: data_out = 8'h9D;
                    16'h4A54: data_out = 8'h9E;
                    16'h4A55: data_out = 8'h9F;
                    16'h4A56: data_out = 8'hA0;
                    16'h4A57: data_out = 8'hA1;
                    16'h4A58: data_out = 8'hA2;
                    16'h4A59: data_out = 8'hA3;
                    16'h4A5A: data_out = 8'hA4;
                    16'h4A5B: data_out = 8'hA5;
                    16'h4A5C: data_out = 8'hA6;
                    16'h4A5D: data_out = 8'hA7;
                    16'h4A5E: data_out = 8'hA8;
                    16'h4A5F: data_out = 8'hA9;
                    16'h4A60: data_out = 8'hAA;
                    16'h4A61: data_out = 8'hAB;
                    16'h4A62: data_out = 8'hAC;
                    16'h4A63: data_out = 8'hAD;
                    16'h4A64: data_out = 8'hAE;
                    16'h4A65: data_out = 8'hAF;
                    16'h4A66: data_out = 8'hB0;
                    16'h4A67: data_out = 8'hB1;
                    16'h4A68: data_out = 8'hB2;
                    16'h4A69: data_out = 8'hB3;
                    16'h4A6A: data_out = 8'hB4;
                    16'h4A6B: data_out = 8'hB5;
                    16'h4A6C: data_out = 8'hB6;
                    16'h4A6D: data_out = 8'hB7;
                    16'h4A6E: data_out = 8'hB8;
                    16'h4A6F: data_out = 8'hB9;
                    16'h4A70: data_out = 8'hBA;
                    16'h4A71: data_out = 8'hBB;
                    16'h4A72: data_out = 8'hBC;
                    16'h4A73: data_out = 8'hBD;
                    16'h4A74: data_out = 8'hBE;
                    16'h4A75: data_out = 8'hBF;
                    16'h4A76: data_out = 8'hC0;
                    16'h4A77: data_out = 8'hC1;
                    16'h4A78: data_out = 8'hC2;
                    16'h4A79: data_out = 8'hC3;
                    16'h4A7A: data_out = 8'hC4;
                    16'h4A7B: data_out = 8'hC5;
                    16'h4A7C: data_out = 8'hC6;
                    16'h4A7D: data_out = 8'hC7;
                    16'h4A7E: data_out = 8'hC8;
                    16'h4A7F: data_out = 8'hC9;
                    16'h4A80: data_out = 8'h4A;
                    16'h4A81: data_out = 8'h49;
                    16'h4A82: data_out = 8'h48;
                    16'h4A83: data_out = 8'h47;
                    16'h4A84: data_out = 8'h46;
                    16'h4A85: data_out = 8'h45;
                    16'h4A86: data_out = 8'h44;
                    16'h4A87: data_out = 8'h43;
                    16'h4A88: data_out = 8'h42;
                    16'h4A89: data_out = 8'h41;
                    16'h4A8A: data_out = 8'h40;
                    16'h4A8B: data_out = 8'h3F;
                    16'h4A8C: data_out = 8'h3E;
                    16'h4A8D: data_out = 8'h3D;
                    16'h4A8E: data_out = 8'h3C;
                    16'h4A8F: data_out = 8'h3B;
                    16'h4A90: data_out = 8'h3A;
                    16'h4A91: data_out = 8'h39;
                    16'h4A92: data_out = 8'h38;
                    16'h4A93: data_out = 8'h37;
                    16'h4A94: data_out = 8'h36;
                    16'h4A95: data_out = 8'h35;
                    16'h4A96: data_out = 8'h34;
                    16'h4A97: data_out = 8'h33;
                    16'h4A98: data_out = 8'h32;
                    16'h4A99: data_out = 8'h31;
                    16'h4A9A: data_out = 8'h30;
                    16'h4A9B: data_out = 8'h2F;
                    16'h4A9C: data_out = 8'h2E;
                    16'h4A9D: data_out = 8'h2D;
                    16'h4A9E: data_out = 8'h2C;
                    16'h4A9F: data_out = 8'h2B;
                    16'h4AA0: data_out = 8'h2A;
                    16'h4AA1: data_out = 8'h29;
                    16'h4AA2: data_out = 8'h28;
                    16'h4AA3: data_out = 8'h27;
                    16'h4AA4: data_out = 8'h26;
                    16'h4AA5: data_out = 8'h25;
                    16'h4AA6: data_out = 8'h24;
                    16'h4AA7: data_out = 8'h23;
                    16'h4AA8: data_out = 8'h22;
                    16'h4AA9: data_out = 8'h21;
                    16'h4AAA: data_out = 8'h20;
                    16'h4AAB: data_out = 8'h1F;
                    16'h4AAC: data_out = 8'h1E;
                    16'h4AAD: data_out = 8'h1D;
                    16'h4AAE: data_out = 8'h1C;
                    16'h4AAF: data_out = 8'h1B;
                    16'h4AB0: data_out = 8'h1A;
                    16'h4AB1: data_out = 8'h19;
                    16'h4AB2: data_out = 8'h18;
                    16'h4AB3: data_out = 8'h17;
                    16'h4AB4: data_out = 8'h16;
                    16'h4AB5: data_out = 8'h15;
                    16'h4AB6: data_out = 8'h14;
                    16'h4AB7: data_out = 8'h13;
                    16'h4AB8: data_out = 8'h12;
                    16'h4AB9: data_out = 8'h11;
                    16'h4ABA: data_out = 8'h10;
                    16'h4ABB: data_out = 8'hF;
                    16'h4ABC: data_out = 8'hE;
                    16'h4ABD: data_out = 8'hD;
                    16'h4ABE: data_out = 8'hC;
                    16'h4ABF: data_out = 8'hB;
                    16'h4AC0: data_out = 8'hA;
                    16'h4AC1: data_out = 8'h9;
                    16'h4AC2: data_out = 8'h8;
                    16'h4AC3: data_out = 8'h7;
                    16'h4AC4: data_out = 8'h6;
                    16'h4AC5: data_out = 8'h5;
                    16'h4AC6: data_out = 8'h4;
                    16'h4AC7: data_out = 8'h3;
                    16'h4AC8: data_out = 8'h2;
                    16'h4AC9: data_out = 8'h1;
                    16'h4ACA: data_out = 8'h0;
                    16'h4ACB: data_out = 8'h81;
                    16'h4ACC: data_out = 8'h82;
                    16'h4ACD: data_out = 8'h83;
                    16'h4ACE: data_out = 8'h84;
                    16'h4ACF: data_out = 8'h85;
                    16'h4AD0: data_out = 8'h86;
                    16'h4AD1: data_out = 8'h87;
                    16'h4AD2: data_out = 8'h88;
                    16'h4AD3: data_out = 8'h89;
                    16'h4AD4: data_out = 8'h8A;
                    16'h4AD5: data_out = 8'h8B;
                    16'h4AD6: data_out = 8'h8C;
                    16'h4AD7: data_out = 8'h8D;
                    16'h4AD8: data_out = 8'h8E;
                    16'h4AD9: data_out = 8'h8F;
                    16'h4ADA: data_out = 8'h90;
                    16'h4ADB: data_out = 8'h91;
                    16'h4ADC: data_out = 8'h92;
                    16'h4ADD: data_out = 8'h93;
                    16'h4ADE: data_out = 8'h94;
                    16'h4ADF: data_out = 8'h95;
                    16'h4AE0: data_out = 8'h96;
                    16'h4AE1: data_out = 8'h97;
                    16'h4AE2: data_out = 8'h98;
                    16'h4AE3: data_out = 8'h99;
                    16'h4AE4: data_out = 8'h9A;
                    16'h4AE5: data_out = 8'h9B;
                    16'h4AE6: data_out = 8'h9C;
                    16'h4AE7: data_out = 8'h9D;
                    16'h4AE8: data_out = 8'h9E;
                    16'h4AE9: data_out = 8'h9F;
                    16'h4AEA: data_out = 8'hA0;
                    16'h4AEB: data_out = 8'hA1;
                    16'h4AEC: data_out = 8'hA2;
                    16'h4AED: data_out = 8'hA3;
                    16'h4AEE: data_out = 8'hA4;
                    16'h4AEF: data_out = 8'hA5;
                    16'h4AF0: data_out = 8'hA6;
                    16'h4AF1: data_out = 8'hA7;
                    16'h4AF2: data_out = 8'hA8;
                    16'h4AF3: data_out = 8'hA9;
                    16'h4AF4: data_out = 8'hAA;
                    16'h4AF5: data_out = 8'hAB;
                    16'h4AF6: data_out = 8'hAC;
                    16'h4AF7: data_out = 8'hAD;
                    16'h4AF8: data_out = 8'hAE;
                    16'h4AF9: data_out = 8'hAF;
                    16'h4AFA: data_out = 8'hB0;
                    16'h4AFB: data_out = 8'hB1;
                    16'h4AFC: data_out = 8'hB2;
                    16'h4AFD: data_out = 8'hB3;
                    16'h4AFE: data_out = 8'hB4;
                    16'h4AFF: data_out = 8'hB5;
                    16'h4B00: data_out = 8'h4B;
                    16'h4B01: data_out = 8'h4C;
                    16'h4B02: data_out = 8'h4D;
                    16'h4B03: data_out = 8'h4E;
                    16'h4B04: data_out = 8'h4F;
                    16'h4B05: data_out = 8'h50;
                    16'h4B06: data_out = 8'h51;
                    16'h4B07: data_out = 8'h52;
                    16'h4B08: data_out = 8'h53;
                    16'h4B09: data_out = 8'h54;
                    16'h4B0A: data_out = 8'h55;
                    16'h4B0B: data_out = 8'h56;
                    16'h4B0C: data_out = 8'h57;
                    16'h4B0D: data_out = 8'h58;
                    16'h4B0E: data_out = 8'h59;
                    16'h4B0F: data_out = 8'h5A;
                    16'h4B10: data_out = 8'h5B;
                    16'h4B11: data_out = 8'h5C;
                    16'h4B12: data_out = 8'h5D;
                    16'h4B13: data_out = 8'h5E;
                    16'h4B14: data_out = 8'h5F;
                    16'h4B15: data_out = 8'h60;
                    16'h4B16: data_out = 8'h61;
                    16'h4B17: data_out = 8'h62;
                    16'h4B18: data_out = 8'h63;
                    16'h4B19: data_out = 8'h64;
                    16'h4B1A: data_out = 8'h65;
                    16'h4B1B: data_out = 8'h66;
                    16'h4B1C: data_out = 8'h67;
                    16'h4B1D: data_out = 8'h68;
                    16'h4B1E: data_out = 8'h69;
                    16'h4B1F: data_out = 8'h6A;
                    16'h4B20: data_out = 8'h6B;
                    16'h4B21: data_out = 8'h6C;
                    16'h4B22: data_out = 8'h6D;
                    16'h4B23: data_out = 8'h6E;
                    16'h4B24: data_out = 8'h6F;
                    16'h4B25: data_out = 8'h70;
                    16'h4B26: data_out = 8'h71;
                    16'h4B27: data_out = 8'h72;
                    16'h4B28: data_out = 8'h73;
                    16'h4B29: data_out = 8'h74;
                    16'h4B2A: data_out = 8'h75;
                    16'h4B2B: data_out = 8'h76;
                    16'h4B2C: data_out = 8'h77;
                    16'h4B2D: data_out = 8'h78;
                    16'h4B2E: data_out = 8'h79;
                    16'h4B2F: data_out = 8'h7A;
                    16'h4B30: data_out = 8'h7B;
                    16'h4B31: data_out = 8'h7C;
                    16'h4B32: data_out = 8'h7D;
                    16'h4B33: data_out = 8'h7E;
                    16'h4B34: data_out = 8'h7F;
                    16'h4B35: data_out = 8'h80;
                    16'h4B36: data_out = 8'h81;
                    16'h4B37: data_out = 8'h82;
                    16'h4B38: data_out = 8'h83;
                    16'h4B39: data_out = 8'h84;
                    16'h4B3A: data_out = 8'h85;
                    16'h4B3B: data_out = 8'h86;
                    16'h4B3C: data_out = 8'h87;
                    16'h4B3D: data_out = 8'h88;
                    16'h4B3E: data_out = 8'h89;
                    16'h4B3F: data_out = 8'h8A;
                    16'h4B40: data_out = 8'h8B;
                    16'h4B41: data_out = 8'h8C;
                    16'h4B42: data_out = 8'h8D;
                    16'h4B43: data_out = 8'h8E;
                    16'h4B44: data_out = 8'h8F;
                    16'h4B45: data_out = 8'h90;
                    16'h4B46: data_out = 8'h91;
                    16'h4B47: data_out = 8'h92;
                    16'h4B48: data_out = 8'h93;
                    16'h4B49: data_out = 8'h94;
                    16'h4B4A: data_out = 8'h95;
                    16'h4B4B: data_out = 8'h96;
                    16'h4B4C: data_out = 8'h97;
                    16'h4B4D: data_out = 8'h98;
                    16'h4B4E: data_out = 8'h99;
                    16'h4B4F: data_out = 8'h9A;
                    16'h4B50: data_out = 8'h9B;
                    16'h4B51: data_out = 8'h9C;
                    16'h4B52: data_out = 8'h9D;
                    16'h4B53: data_out = 8'h9E;
                    16'h4B54: data_out = 8'h9F;
                    16'h4B55: data_out = 8'hA0;
                    16'h4B56: data_out = 8'hA1;
                    16'h4B57: data_out = 8'hA2;
                    16'h4B58: data_out = 8'hA3;
                    16'h4B59: data_out = 8'hA4;
                    16'h4B5A: data_out = 8'hA5;
                    16'h4B5B: data_out = 8'hA6;
                    16'h4B5C: data_out = 8'hA7;
                    16'h4B5D: data_out = 8'hA8;
                    16'h4B5E: data_out = 8'hA9;
                    16'h4B5F: data_out = 8'hAA;
                    16'h4B60: data_out = 8'hAB;
                    16'h4B61: data_out = 8'hAC;
                    16'h4B62: data_out = 8'hAD;
                    16'h4B63: data_out = 8'hAE;
                    16'h4B64: data_out = 8'hAF;
                    16'h4B65: data_out = 8'hB0;
                    16'h4B66: data_out = 8'hB1;
                    16'h4B67: data_out = 8'hB2;
                    16'h4B68: data_out = 8'hB3;
                    16'h4B69: data_out = 8'hB4;
                    16'h4B6A: data_out = 8'hB5;
                    16'h4B6B: data_out = 8'hB6;
                    16'h4B6C: data_out = 8'hB7;
                    16'h4B6D: data_out = 8'hB8;
                    16'h4B6E: data_out = 8'hB9;
                    16'h4B6F: data_out = 8'hBA;
                    16'h4B70: data_out = 8'hBB;
                    16'h4B71: data_out = 8'hBC;
                    16'h4B72: data_out = 8'hBD;
                    16'h4B73: data_out = 8'hBE;
                    16'h4B74: data_out = 8'hBF;
                    16'h4B75: data_out = 8'hC0;
                    16'h4B76: data_out = 8'hC1;
                    16'h4B77: data_out = 8'hC2;
                    16'h4B78: data_out = 8'hC3;
                    16'h4B79: data_out = 8'hC4;
                    16'h4B7A: data_out = 8'hC5;
                    16'h4B7B: data_out = 8'hC6;
                    16'h4B7C: data_out = 8'hC7;
                    16'h4B7D: data_out = 8'hC8;
                    16'h4B7E: data_out = 8'hC9;
                    16'h4B7F: data_out = 8'hCA;
                    16'h4B80: data_out = 8'h4B;
                    16'h4B81: data_out = 8'h4A;
                    16'h4B82: data_out = 8'h49;
                    16'h4B83: data_out = 8'h48;
                    16'h4B84: data_out = 8'h47;
                    16'h4B85: data_out = 8'h46;
                    16'h4B86: data_out = 8'h45;
                    16'h4B87: data_out = 8'h44;
                    16'h4B88: data_out = 8'h43;
                    16'h4B89: data_out = 8'h42;
                    16'h4B8A: data_out = 8'h41;
                    16'h4B8B: data_out = 8'h40;
                    16'h4B8C: data_out = 8'h3F;
                    16'h4B8D: data_out = 8'h3E;
                    16'h4B8E: data_out = 8'h3D;
                    16'h4B8F: data_out = 8'h3C;
                    16'h4B90: data_out = 8'h3B;
                    16'h4B91: data_out = 8'h3A;
                    16'h4B92: data_out = 8'h39;
                    16'h4B93: data_out = 8'h38;
                    16'h4B94: data_out = 8'h37;
                    16'h4B95: data_out = 8'h36;
                    16'h4B96: data_out = 8'h35;
                    16'h4B97: data_out = 8'h34;
                    16'h4B98: data_out = 8'h33;
                    16'h4B99: data_out = 8'h32;
                    16'h4B9A: data_out = 8'h31;
                    16'h4B9B: data_out = 8'h30;
                    16'h4B9C: data_out = 8'h2F;
                    16'h4B9D: data_out = 8'h2E;
                    16'h4B9E: data_out = 8'h2D;
                    16'h4B9F: data_out = 8'h2C;
                    16'h4BA0: data_out = 8'h2B;
                    16'h4BA1: data_out = 8'h2A;
                    16'h4BA2: data_out = 8'h29;
                    16'h4BA3: data_out = 8'h28;
                    16'h4BA4: data_out = 8'h27;
                    16'h4BA5: data_out = 8'h26;
                    16'h4BA6: data_out = 8'h25;
                    16'h4BA7: data_out = 8'h24;
                    16'h4BA8: data_out = 8'h23;
                    16'h4BA9: data_out = 8'h22;
                    16'h4BAA: data_out = 8'h21;
                    16'h4BAB: data_out = 8'h20;
                    16'h4BAC: data_out = 8'h1F;
                    16'h4BAD: data_out = 8'h1E;
                    16'h4BAE: data_out = 8'h1D;
                    16'h4BAF: data_out = 8'h1C;
                    16'h4BB0: data_out = 8'h1B;
                    16'h4BB1: data_out = 8'h1A;
                    16'h4BB2: data_out = 8'h19;
                    16'h4BB3: data_out = 8'h18;
                    16'h4BB4: data_out = 8'h17;
                    16'h4BB5: data_out = 8'h16;
                    16'h4BB6: data_out = 8'h15;
                    16'h4BB7: data_out = 8'h14;
                    16'h4BB8: data_out = 8'h13;
                    16'h4BB9: data_out = 8'h12;
                    16'h4BBA: data_out = 8'h11;
                    16'h4BBB: data_out = 8'h10;
                    16'h4BBC: data_out = 8'hF;
                    16'h4BBD: data_out = 8'hE;
                    16'h4BBE: data_out = 8'hD;
                    16'h4BBF: data_out = 8'hC;
                    16'h4BC0: data_out = 8'hB;
                    16'h4BC1: data_out = 8'hA;
                    16'h4BC2: data_out = 8'h9;
                    16'h4BC3: data_out = 8'h8;
                    16'h4BC4: data_out = 8'h7;
                    16'h4BC5: data_out = 8'h6;
                    16'h4BC6: data_out = 8'h5;
                    16'h4BC7: data_out = 8'h4;
                    16'h4BC8: data_out = 8'h3;
                    16'h4BC9: data_out = 8'h2;
                    16'h4BCA: data_out = 8'h1;
                    16'h4BCB: data_out = 8'h0;
                    16'h4BCC: data_out = 8'h81;
                    16'h4BCD: data_out = 8'h82;
                    16'h4BCE: data_out = 8'h83;
                    16'h4BCF: data_out = 8'h84;
                    16'h4BD0: data_out = 8'h85;
                    16'h4BD1: data_out = 8'h86;
                    16'h4BD2: data_out = 8'h87;
                    16'h4BD3: data_out = 8'h88;
                    16'h4BD4: data_out = 8'h89;
                    16'h4BD5: data_out = 8'h8A;
                    16'h4BD6: data_out = 8'h8B;
                    16'h4BD7: data_out = 8'h8C;
                    16'h4BD8: data_out = 8'h8D;
                    16'h4BD9: data_out = 8'h8E;
                    16'h4BDA: data_out = 8'h8F;
                    16'h4BDB: data_out = 8'h90;
                    16'h4BDC: data_out = 8'h91;
                    16'h4BDD: data_out = 8'h92;
                    16'h4BDE: data_out = 8'h93;
                    16'h4BDF: data_out = 8'h94;
                    16'h4BE0: data_out = 8'h95;
                    16'h4BE1: data_out = 8'h96;
                    16'h4BE2: data_out = 8'h97;
                    16'h4BE3: data_out = 8'h98;
                    16'h4BE4: data_out = 8'h99;
                    16'h4BE5: data_out = 8'h9A;
                    16'h4BE6: data_out = 8'h9B;
                    16'h4BE7: data_out = 8'h9C;
                    16'h4BE8: data_out = 8'h9D;
                    16'h4BE9: data_out = 8'h9E;
                    16'h4BEA: data_out = 8'h9F;
                    16'h4BEB: data_out = 8'hA0;
                    16'h4BEC: data_out = 8'hA1;
                    16'h4BED: data_out = 8'hA2;
                    16'h4BEE: data_out = 8'hA3;
                    16'h4BEF: data_out = 8'hA4;
                    16'h4BF0: data_out = 8'hA5;
                    16'h4BF1: data_out = 8'hA6;
                    16'h4BF2: data_out = 8'hA7;
                    16'h4BF3: data_out = 8'hA8;
                    16'h4BF4: data_out = 8'hA9;
                    16'h4BF5: data_out = 8'hAA;
                    16'h4BF6: data_out = 8'hAB;
                    16'h4BF7: data_out = 8'hAC;
                    16'h4BF8: data_out = 8'hAD;
                    16'h4BF9: data_out = 8'hAE;
                    16'h4BFA: data_out = 8'hAF;
                    16'h4BFB: data_out = 8'hB0;
                    16'h4BFC: data_out = 8'hB1;
                    16'h4BFD: data_out = 8'hB2;
                    16'h4BFE: data_out = 8'hB3;
                    16'h4BFF: data_out = 8'hB4;
                    16'h4C00: data_out = 8'h4C;
                    16'h4C01: data_out = 8'h4D;
                    16'h4C02: data_out = 8'h4E;
                    16'h4C03: data_out = 8'h4F;
                    16'h4C04: data_out = 8'h50;
                    16'h4C05: data_out = 8'h51;
                    16'h4C06: data_out = 8'h52;
                    16'h4C07: data_out = 8'h53;
                    16'h4C08: data_out = 8'h54;
                    16'h4C09: data_out = 8'h55;
                    16'h4C0A: data_out = 8'h56;
                    16'h4C0B: data_out = 8'h57;
                    16'h4C0C: data_out = 8'h58;
                    16'h4C0D: data_out = 8'h59;
                    16'h4C0E: data_out = 8'h5A;
                    16'h4C0F: data_out = 8'h5B;
                    16'h4C10: data_out = 8'h5C;
                    16'h4C11: data_out = 8'h5D;
                    16'h4C12: data_out = 8'h5E;
                    16'h4C13: data_out = 8'h5F;
                    16'h4C14: data_out = 8'h60;
                    16'h4C15: data_out = 8'h61;
                    16'h4C16: data_out = 8'h62;
                    16'h4C17: data_out = 8'h63;
                    16'h4C18: data_out = 8'h64;
                    16'h4C19: data_out = 8'h65;
                    16'h4C1A: data_out = 8'h66;
                    16'h4C1B: data_out = 8'h67;
                    16'h4C1C: data_out = 8'h68;
                    16'h4C1D: data_out = 8'h69;
                    16'h4C1E: data_out = 8'h6A;
                    16'h4C1F: data_out = 8'h6B;
                    16'h4C20: data_out = 8'h6C;
                    16'h4C21: data_out = 8'h6D;
                    16'h4C22: data_out = 8'h6E;
                    16'h4C23: data_out = 8'h6F;
                    16'h4C24: data_out = 8'h70;
                    16'h4C25: data_out = 8'h71;
                    16'h4C26: data_out = 8'h72;
                    16'h4C27: data_out = 8'h73;
                    16'h4C28: data_out = 8'h74;
                    16'h4C29: data_out = 8'h75;
                    16'h4C2A: data_out = 8'h76;
                    16'h4C2B: data_out = 8'h77;
                    16'h4C2C: data_out = 8'h78;
                    16'h4C2D: data_out = 8'h79;
                    16'h4C2E: data_out = 8'h7A;
                    16'h4C2F: data_out = 8'h7B;
                    16'h4C30: data_out = 8'h7C;
                    16'h4C31: data_out = 8'h7D;
                    16'h4C32: data_out = 8'h7E;
                    16'h4C33: data_out = 8'h7F;
                    16'h4C34: data_out = 8'h80;
                    16'h4C35: data_out = 8'h81;
                    16'h4C36: data_out = 8'h82;
                    16'h4C37: data_out = 8'h83;
                    16'h4C38: data_out = 8'h84;
                    16'h4C39: data_out = 8'h85;
                    16'h4C3A: data_out = 8'h86;
                    16'h4C3B: data_out = 8'h87;
                    16'h4C3C: data_out = 8'h88;
                    16'h4C3D: data_out = 8'h89;
                    16'h4C3E: data_out = 8'h8A;
                    16'h4C3F: data_out = 8'h8B;
                    16'h4C40: data_out = 8'h8C;
                    16'h4C41: data_out = 8'h8D;
                    16'h4C42: data_out = 8'h8E;
                    16'h4C43: data_out = 8'h8F;
                    16'h4C44: data_out = 8'h90;
                    16'h4C45: data_out = 8'h91;
                    16'h4C46: data_out = 8'h92;
                    16'h4C47: data_out = 8'h93;
                    16'h4C48: data_out = 8'h94;
                    16'h4C49: data_out = 8'h95;
                    16'h4C4A: data_out = 8'h96;
                    16'h4C4B: data_out = 8'h97;
                    16'h4C4C: data_out = 8'h98;
                    16'h4C4D: data_out = 8'h99;
                    16'h4C4E: data_out = 8'h9A;
                    16'h4C4F: data_out = 8'h9B;
                    16'h4C50: data_out = 8'h9C;
                    16'h4C51: data_out = 8'h9D;
                    16'h4C52: data_out = 8'h9E;
                    16'h4C53: data_out = 8'h9F;
                    16'h4C54: data_out = 8'hA0;
                    16'h4C55: data_out = 8'hA1;
                    16'h4C56: data_out = 8'hA2;
                    16'h4C57: data_out = 8'hA3;
                    16'h4C58: data_out = 8'hA4;
                    16'h4C59: data_out = 8'hA5;
                    16'h4C5A: data_out = 8'hA6;
                    16'h4C5B: data_out = 8'hA7;
                    16'h4C5C: data_out = 8'hA8;
                    16'h4C5D: data_out = 8'hA9;
                    16'h4C5E: data_out = 8'hAA;
                    16'h4C5F: data_out = 8'hAB;
                    16'h4C60: data_out = 8'hAC;
                    16'h4C61: data_out = 8'hAD;
                    16'h4C62: data_out = 8'hAE;
                    16'h4C63: data_out = 8'hAF;
                    16'h4C64: data_out = 8'hB0;
                    16'h4C65: data_out = 8'hB1;
                    16'h4C66: data_out = 8'hB2;
                    16'h4C67: data_out = 8'hB3;
                    16'h4C68: data_out = 8'hB4;
                    16'h4C69: data_out = 8'hB5;
                    16'h4C6A: data_out = 8'hB6;
                    16'h4C6B: data_out = 8'hB7;
                    16'h4C6C: data_out = 8'hB8;
                    16'h4C6D: data_out = 8'hB9;
                    16'h4C6E: data_out = 8'hBA;
                    16'h4C6F: data_out = 8'hBB;
                    16'h4C70: data_out = 8'hBC;
                    16'h4C71: data_out = 8'hBD;
                    16'h4C72: data_out = 8'hBE;
                    16'h4C73: data_out = 8'hBF;
                    16'h4C74: data_out = 8'hC0;
                    16'h4C75: data_out = 8'hC1;
                    16'h4C76: data_out = 8'hC2;
                    16'h4C77: data_out = 8'hC3;
                    16'h4C78: data_out = 8'hC4;
                    16'h4C79: data_out = 8'hC5;
                    16'h4C7A: data_out = 8'hC6;
                    16'h4C7B: data_out = 8'hC7;
                    16'h4C7C: data_out = 8'hC8;
                    16'h4C7D: data_out = 8'hC9;
                    16'h4C7E: data_out = 8'hCA;
                    16'h4C7F: data_out = 8'hCB;
                    16'h4C80: data_out = 8'h4C;
                    16'h4C81: data_out = 8'h4B;
                    16'h4C82: data_out = 8'h4A;
                    16'h4C83: data_out = 8'h49;
                    16'h4C84: data_out = 8'h48;
                    16'h4C85: data_out = 8'h47;
                    16'h4C86: data_out = 8'h46;
                    16'h4C87: data_out = 8'h45;
                    16'h4C88: data_out = 8'h44;
                    16'h4C89: data_out = 8'h43;
                    16'h4C8A: data_out = 8'h42;
                    16'h4C8B: data_out = 8'h41;
                    16'h4C8C: data_out = 8'h40;
                    16'h4C8D: data_out = 8'h3F;
                    16'h4C8E: data_out = 8'h3E;
                    16'h4C8F: data_out = 8'h3D;
                    16'h4C90: data_out = 8'h3C;
                    16'h4C91: data_out = 8'h3B;
                    16'h4C92: data_out = 8'h3A;
                    16'h4C93: data_out = 8'h39;
                    16'h4C94: data_out = 8'h38;
                    16'h4C95: data_out = 8'h37;
                    16'h4C96: data_out = 8'h36;
                    16'h4C97: data_out = 8'h35;
                    16'h4C98: data_out = 8'h34;
                    16'h4C99: data_out = 8'h33;
                    16'h4C9A: data_out = 8'h32;
                    16'h4C9B: data_out = 8'h31;
                    16'h4C9C: data_out = 8'h30;
                    16'h4C9D: data_out = 8'h2F;
                    16'h4C9E: data_out = 8'h2E;
                    16'h4C9F: data_out = 8'h2D;
                    16'h4CA0: data_out = 8'h2C;
                    16'h4CA1: data_out = 8'h2B;
                    16'h4CA2: data_out = 8'h2A;
                    16'h4CA3: data_out = 8'h29;
                    16'h4CA4: data_out = 8'h28;
                    16'h4CA5: data_out = 8'h27;
                    16'h4CA6: data_out = 8'h26;
                    16'h4CA7: data_out = 8'h25;
                    16'h4CA8: data_out = 8'h24;
                    16'h4CA9: data_out = 8'h23;
                    16'h4CAA: data_out = 8'h22;
                    16'h4CAB: data_out = 8'h21;
                    16'h4CAC: data_out = 8'h20;
                    16'h4CAD: data_out = 8'h1F;
                    16'h4CAE: data_out = 8'h1E;
                    16'h4CAF: data_out = 8'h1D;
                    16'h4CB0: data_out = 8'h1C;
                    16'h4CB1: data_out = 8'h1B;
                    16'h4CB2: data_out = 8'h1A;
                    16'h4CB3: data_out = 8'h19;
                    16'h4CB4: data_out = 8'h18;
                    16'h4CB5: data_out = 8'h17;
                    16'h4CB6: data_out = 8'h16;
                    16'h4CB7: data_out = 8'h15;
                    16'h4CB8: data_out = 8'h14;
                    16'h4CB9: data_out = 8'h13;
                    16'h4CBA: data_out = 8'h12;
                    16'h4CBB: data_out = 8'h11;
                    16'h4CBC: data_out = 8'h10;
                    16'h4CBD: data_out = 8'hF;
                    16'h4CBE: data_out = 8'hE;
                    16'h4CBF: data_out = 8'hD;
                    16'h4CC0: data_out = 8'hC;
                    16'h4CC1: data_out = 8'hB;
                    16'h4CC2: data_out = 8'hA;
                    16'h4CC3: data_out = 8'h9;
                    16'h4CC4: data_out = 8'h8;
                    16'h4CC5: data_out = 8'h7;
                    16'h4CC6: data_out = 8'h6;
                    16'h4CC7: data_out = 8'h5;
                    16'h4CC8: data_out = 8'h4;
                    16'h4CC9: data_out = 8'h3;
                    16'h4CCA: data_out = 8'h2;
                    16'h4CCB: data_out = 8'h1;
                    16'h4CCC: data_out = 8'h0;
                    16'h4CCD: data_out = 8'h81;
                    16'h4CCE: data_out = 8'h82;
                    16'h4CCF: data_out = 8'h83;
                    16'h4CD0: data_out = 8'h84;
                    16'h4CD1: data_out = 8'h85;
                    16'h4CD2: data_out = 8'h86;
                    16'h4CD3: data_out = 8'h87;
                    16'h4CD4: data_out = 8'h88;
                    16'h4CD5: data_out = 8'h89;
                    16'h4CD6: data_out = 8'h8A;
                    16'h4CD7: data_out = 8'h8B;
                    16'h4CD8: data_out = 8'h8C;
                    16'h4CD9: data_out = 8'h8D;
                    16'h4CDA: data_out = 8'h8E;
                    16'h4CDB: data_out = 8'h8F;
                    16'h4CDC: data_out = 8'h90;
                    16'h4CDD: data_out = 8'h91;
                    16'h4CDE: data_out = 8'h92;
                    16'h4CDF: data_out = 8'h93;
                    16'h4CE0: data_out = 8'h94;
                    16'h4CE1: data_out = 8'h95;
                    16'h4CE2: data_out = 8'h96;
                    16'h4CE3: data_out = 8'h97;
                    16'h4CE4: data_out = 8'h98;
                    16'h4CE5: data_out = 8'h99;
                    16'h4CE6: data_out = 8'h9A;
                    16'h4CE7: data_out = 8'h9B;
                    16'h4CE8: data_out = 8'h9C;
                    16'h4CE9: data_out = 8'h9D;
                    16'h4CEA: data_out = 8'h9E;
                    16'h4CEB: data_out = 8'h9F;
                    16'h4CEC: data_out = 8'hA0;
                    16'h4CED: data_out = 8'hA1;
                    16'h4CEE: data_out = 8'hA2;
                    16'h4CEF: data_out = 8'hA3;
                    16'h4CF0: data_out = 8'hA4;
                    16'h4CF1: data_out = 8'hA5;
                    16'h4CF2: data_out = 8'hA6;
                    16'h4CF3: data_out = 8'hA7;
                    16'h4CF4: data_out = 8'hA8;
                    16'h4CF5: data_out = 8'hA9;
                    16'h4CF6: data_out = 8'hAA;
                    16'h4CF7: data_out = 8'hAB;
                    16'h4CF8: data_out = 8'hAC;
                    16'h4CF9: data_out = 8'hAD;
                    16'h4CFA: data_out = 8'hAE;
                    16'h4CFB: data_out = 8'hAF;
                    16'h4CFC: data_out = 8'hB0;
                    16'h4CFD: data_out = 8'hB1;
                    16'h4CFE: data_out = 8'hB2;
                    16'h4CFF: data_out = 8'hB3;
                    16'h4D00: data_out = 8'h4D;
                    16'h4D01: data_out = 8'h4E;
                    16'h4D02: data_out = 8'h4F;
                    16'h4D03: data_out = 8'h50;
                    16'h4D04: data_out = 8'h51;
                    16'h4D05: data_out = 8'h52;
                    16'h4D06: data_out = 8'h53;
                    16'h4D07: data_out = 8'h54;
                    16'h4D08: data_out = 8'h55;
                    16'h4D09: data_out = 8'h56;
                    16'h4D0A: data_out = 8'h57;
                    16'h4D0B: data_out = 8'h58;
                    16'h4D0C: data_out = 8'h59;
                    16'h4D0D: data_out = 8'h5A;
                    16'h4D0E: data_out = 8'h5B;
                    16'h4D0F: data_out = 8'h5C;
                    16'h4D10: data_out = 8'h5D;
                    16'h4D11: data_out = 8'h5E;
                    16'h4D12: data_out = 8'h5F;
                    16'h4D13: data_out = 8'h60;
                    16'h4D14: data_out = 8'h61;
                    16'h4D15: data_out = 8'h62;
                    16'h4D16: data_out = 8'h63;
                    16'h4D17: data_out = 8'h64;
                    16'h4D18: data_out = 8'h65;
                    16'h4D19: data_out = 8'h66;
                    16'h4D1A: data_out = 8'h67;
                    16'h4D1B: data_out = 8'h68;
                    16'h4D1C: data_out = 8'h69;
                    16'h4D1D: data_out = 8'h6A;
                    16'h4D1E: data_out = 8'h6B;
                    16'h4D1F: data_out = 8'h6C;
                    16'h4D20: data_out = 8'h6D;
                    16'h4D21: data_out = 8'h6E;
                    16'h4D22: data_out = 8'h6F;
                    16'h4D23: data_out = 8'h70;
                    16'h4D24: data_out = 8'h71;
                    16'h4D25: data_out = 8'h72;
                    16'h4D26: data_out = 8'h73;
                    16'h4D27: data_out = 8'h74;
                    16'h4D28: data_out = 8'h75;
                    16'h4D29: data_out = 8'h76;
                    16'h4D2A: data_out = 8'h77;
                    16'h4D2B: data_out = 8'h78;
                    16'h4D2C: data_out = 8'h79;
                    16'h4D2D: data_out = 8'h7A;
                    16'h4D2E: data_out = 8'h7B;
                    16'h4D2F: data_out = 8'h7C;
                    16'h4D30: data_out = 8'h7D;
                    16'h4D31: data_out = 8'h7E;
                    16'h4D32: data_out = 8'h7F;
                    16'h4D33: data_out = 8'h80;
                    16'h4D34: data_out = 8'h81;
                    16'h4D35: data_out = 8'h82;
                    16'h4D36: data_out = 8'h83;
                    16'h4D37: data_out = 8'h84;
                    16'h4D38: data_out = 8'h85;
                    16'h4D39: data_out = 8'h86;
                    16'h4D3A: data_out = 8'h87;
                    16'h4D3B: data_out = 8'h88;
                    16'h4D3C: data_out = 8'h89;
                    16'h4D3D: data_out = 8'h8A;
                    16'h4D3E: data_out = 8'h8B;
                    16'h4D3F: data_out = 8'h8C;
                    16'h4D40: data_out = 8'h8D;
                    16'h4D41: data_out = 8'h8E;
                    16'h4D42: data_out = 8'h8F;
                    16'h4D43: data_out = 8'h90;
                    16'h4D44: data_out = 8'h91;
                    16'h4D45: data_out = 8'h92;
                    16'h4D46: data_out = 8'h93;
                    16'h4D47: data_out = 8'h94;
                    16'h4D48: data_out = 8'h95;
                    16'h4D49: data_out = 8'h96;
                    16'h4D4A: data_out = 8'h97;
                    16'h4D4B: data_out = 8'h98;
                    16'h4D4C: data_out = 8'h99;
                    16'h4D4D: data_out = 8'h9A;
                    16'h4D4E: data_out = 8'h9B;
                    16'h4D4F: data_out = 8'h9C;
                    16'h4D50: data_out = 8'h9D;
                    16'h4D51: data_out = 8'h9E;
                    16'h4D52: data_out = 8'h9F;
                    16'h4D53: data_out = 8'hA0;
                    16'h4D54: data_out = 8'hA1;
                    16'h4D55: data_out = 8'hA2;
                    16'h4D56: data_out = 8'hA3;
                    16'h4D57: data_out = 8'hA4;
                    16'h4D58: data_out = 8'hA5;
                    16'h4D59: data_out = 8'hA6;
                    16'h4D5A: data_out = 8'hA7;
                    16'h4D5B: data_out = 8'hA8;
                    16'h4D5C: data_out = 8'hA9;
                    16'h4D5D: data_out = 8'hAA;
                    16'h4D5E: data_out = 8'hAB;
                    16'h4D5F: data_out = 8'hAC;
                    16'h4D60: data_out = 8'hAD;
                    16'h4D61: data_out = 8'hAE;
                    16'h4D62: data_out = 8'hAF;
                    16'h4D63: data_out = 8'hB0;
                    16'h4D64: data_out = 8'hB1;
                    16'h4D65: data_out = 8'hB2;
                    16'h4D66: data_out = 8'hB3;
                    16'h4D67: data_out = 8'hB4;
                    16'h4D68: data_out = 8'hB5;
                    16'h4D69: data_out = 8'hB6;
                    16'h4D6A: data_out = 8'hB7;
                    16'h4D6B: data_out = 8'hB8;
                    16'h4D6C: data_out = 8'hB9;
                    16'h4D6D: data_out = 8'hBA;
                    16'h4D6E: data_out = 8'hBB;
                    16'h4D6F: data_out = 8'hBC;
                    16'h4D70: data_out = 8'hBD;
                    16'h4D71: data_out = 8'hBE;
                    16'h4D72: data_out = 8'hBF;
                    16'h4D73: data_out = 8'hC0;
                    16'h4D74: data_out = 8'hC1;
                    16'h4D75: data_out = 8'hC2;
                    16'h4D76: data_out = 8'hC3;
                    16'h4D77: data_out = 8'hC4;
                    16'h4D78: data_out = 8'hC5;
                    16'h4D79: data_out = 8'hC6;
                    16'h4D7A: data_out = 8'hC7;
                    16'h4D7B: data_out = 8'hC8;
                    16'h4D7C: data_out = 8'hC9;
                    16'h4D7D: data_out = 8'hCA;
                    16'h4D7E: data_out = 8'hCB;
                    16'h4D7F: data_out = 8'hCC;
                    16'h4D80: data_out = 8'h4D;
                    16'h4D81: data_out = 8'h4C;
                    16'h4D82: data_out = 8'h4B;
                    16'h4D83: data_out = 8'h4A;
                    16'h4D84: data_out = 8'h49;
                    16'h4D85: data_out = 8'h48;
                    16'h4D86: data_out = 8'h47;
                    16'h4D87: data_out = 8'h46;
                    16'h4D88: data_out = 8'h45;
                    16'h4D89: data_out = 8'h44;
                    16'h4D8A: data_out = 8'h43;
                    16'h4D8B: data_out = 8'h42;
                    16'h4D8C: data_out = 8'h41;
                    16'h4D8D: data_out = 8'h40;
                    16'h4D8E: data_out = 8'h3F;
                    16'h4D8F: data_out = 8'h3E;
                    16'h4D90: data_out = 8'h3D;
                    16'h4D91: data_out = 8'h3C;
                    16'h4D92: data_out = 8'h3B;
                    16'h4D93: data_out = 8'h3A;
                    16'h4D94: data_out = 8'h39;
                    16'h4D95: data_out = 8'h38;
                    16'h4D96: data_out = 8'h37;
                    16'h4D97: data_out = 8'h36;
                    16'h4D98: data_out = 8'h35;
                    16'h4D99: data_out = 8'h34;
                    16'h4D9A: data_out = 8'h33;
                    16'h4D9B: data_out = 8'h32;
                    16'h4D9C: data_out = 8'h31;
                    16'h4D9D: data_out = 8'h30;
                    16'h4D9E: data_out = 8'h2F;
                    16'h4D9F: data_out = 8'h2E;
                    16'h4DA0: data_out = 8'h2D;
                    16'h4DA1: data_out = 8'h2C;
                    16'h4DA2: data_out = 8'h2B;
                    16'h4DA3: data_out = 8'h2A;
                    16'h4DA4: data_out = 8'h29;
                    16'h4DA5: data_out = 8'h28;
                    16'h4DA6: data_out = 8'h27;
                    16'h4DA7: data_out = 8'h26;
                    16'h4DA8: data_out = 8'h25;
                    16'h4DA9: data_out = 8'h24;
                    16'h4DAA: data_out = 8'h23;
                    16'h4DAB: data_out = 8'h22;
                    16'h4DAC: data_out = 8'h21;
                    16'h4DAD: data_out = 8'h20;
                    16'h4DAE: data_out = 8'h1F;
                    16'h4DAF: data_out = 8'h1E;
                    16'h4DB0: data_out = 8'h1D;
                    16'h4DB1: data_out = 8'h1C;
                    16'h4DB2: data_out = 8'h1B;
                    16'h4DB3: data_out = 8'h1A;
                    16'h4DB4: data_out = 8'h19;
                    16'h4DB5: data_out = 8'h18;
                    16'h4DB6: data_out = 8'h17;
                    16'h4DB7: data_out = 8'h16;
                    16'h4DB8: data_out = 8'h15;
                    16'h4DB9: data_out = 8'h14;
                    16'h4DBA: data_out = 8'h13;
                    16'h4DBB: data_out = 8'h12;
                    16'h4DBC: data_out = 8'h11;
                    16'h4DBD: data_out = 8'h10;
                    16'h4DBE: data_out = 8'hF;
                    16'h4DBF: data_out = 8'hE;
                    16'h4DC0: data_out = 8'hD;
                    16'h4DC1: data_out = 8'hC;
                    16'h4DC2: data_out = 8'hB;
                    16'h4DC3: data_out = 8'hA;
                    16'h4DC4: data_out = 8'h9;
                    16'h4DC5: data_out = 8'h8;
                    16'h4DC6: data_out = 8'h7;
                    16'h4DC7: data_out = 8'h6;
                    16'h4DC8: data_out = 8'h5;
                    16'h4DC9: data_out = 8'h4;
                    16'h4DCA: data_out = 8'h3;
                    16'h4DCB: data_out = 8'h2;
                    16'h4DCC: data_out = 8'h1;
                    16'h4DCD: data_out = 8'h0;
                    16'h4DCE: data_out = 8'h81;
                    16'h4DCF: data_out = 8'h82;
                    16'h4DD0: data_out = 8'h83;
                    16'h4DD1: data_out = 8'h84;
                    16'h4DD2: data_out = 8'h85;
                    16'h4DD3: data_out = 8'h86;
                    16'h4DD4: data_out = 8'h87;
                    16'h4DD5: data_out = 8'h88;
                    16'h4DD6: data_out = 8'h89;
                    16'h4DD7: data_out = 8'h8A;
                    16'h4DD8: data_out = 8'h8B;
                    16'h4DD9: data_out = 8'h8C;
                    16'h4DDA: data_out = 8'h8D;
                    16'h4DDB: data_out = 8'h8E;
                    16'h4DDC: data_out = 8'h8F;
                    16'h4DDD: data_out = 8'h90;
                    16'h4DDE: data_out = 8'h91;
                    16'h4DDF: data_out = 8'h92;
                    16'h4DE0: data_out = 8'h93;
                    16'h4DE1: data_out = 8'h94;
                    16'h4DE2: data_out = 8'h95;
                    16'h4DE3: data_out = 8'h96;
                    16'h4DE4: data_out = 8'h97;
                    16'h4DE5: data_out = 8'h98;
                    16'h4DE6: data_out = 8'h99;
                    16'h4DE7: data_out = 8'h9A;
                    16'h4DE8: data_out = 8'h9B;
                    16'h4DE9: data_out = 8'h9C;
                    16'h4DEA: data_out = 8'h9D;
                    16'h4DEB: data_out = 8'h9E;
                    16'h4DEC: data_out = 8'h9F;
                    16'h4DED: data_out = 8'hA0;
                    16'h4DEE: data_out = 8'hA1;
                    16'h4DEF: data_out = 8'hA2;
                    16'h4DF0: data_out = 8'hA3;
                    16'h4DF1: data_out = 8'hA4;
                    16'h4DF2: data_out = 8'hA5;
                    16'h4DF3: data_out = 8'hA6;
                    16'h4DF4: data_out = 8'hA7;
                    16'h4DF5: data_out = 8'hA8;
                    16'h4DF6: data_out = 8'hA9;
                    16'h4DF7: data_out = 8'hAA;
                    16'h4DF8: data_out = 8'hAB;
                    16'h4DF9: data_out = 8'hAC;
                    16'h4DFA: data_out = 8'hAD;
                    16'h4DFB: data_out = 8'hAE;
                    16'h4DFC: data_out = 8'hAF;
                    16'h4DFD: data_out = 8'hB0;
                    16'h4DFE: data_out = 8'hB1;
                    16'h4DFF: data_out = 8'hB2;
                    16'h4E00: data_out = 8'h4E;
                    16'h4E01: data_out = 8'h4F;
                    16'h4E02: data_out = 8'h50;
                    16'h4E03: data_out = 8'h51;
                    16'h4E04: data_out = 8'h52;
                    16'h4E05: data_out = 8'h53;
                    16'h4E06: data_out = 8'h54;
                    16'h4E07: data_out = 8'h55;
                    16'h4E08: data_out = 8'h56;
                    16'h4E09: data_out = 8'h57;
                    16'h4E0A: data_out = 8'h58;
                    16'h4E0B: data_out = 8'h59;
                    16'h4E0C: data_out = 8'h5A;
                    16'h4E0D: data_out = 8'h5B;
                    16'h4E0E: data_out = 8'h5C;
                    16'h4E0F: data_out = 8'h5D;
                    16'h4E10: data_out = 8'h5E;
                    16'h4E11: data_out = 8'h5F;
                    16'h4E12: data_out = 8'h60;
                    16'h4E13: data_out = 8'h61;
                    16'h4E14: data_out = 8'h62;
                    16'h4E15: data_out = 8'h63;
                    16'h4E16: data_out = 8'h64;
                    16'h4E17: data_out = 8'h65;
                    16'h4E18: data_out = 8'h66;
                    16'h4E19: data_out = 8'h67;
                    16'h4E1A: data_out = 8'h68;
                    16'h4E1B: data_out = 8'h69;
                    16'h4E1C: data_out = 8'h6A;
                    16'h4E1D: data_out = 8'h6B;
                    16'h4E1E: data_out = 8'h6C;
                    16'h4E1F: data_out = 8'h6D;
                    16'h4E20: data_out = 8'h6E;
                    16'h4E21: data_out = 8'h6F;
                    16'h4E22: data_out = 8'h70;
                    16'h4E23: data_out = 8'h71;
                    16'h4E24: data_out = 8'h72;
                    16'h4E25: data_out = 8'h73;
                    16'h4E26: data_out = 8'h74;
                    16'h4E27: data_out = 8'h75;
                    16'h4E28: data_out = 8'h76;
                    16'h4E29: data_out = 8'h77;
                    16'h4E2A: data_out = 8'h78;
                    16'h4E2B: data_out = 8'h79;
                    16'h4E2C: data_out = 8'h7A;
                    16'h4E2D: data_out = 8'h7B;
                    16'h4E2E: data_out = 8'h7C;
                    16'h4E2F: data_out = 8'h7D;
                    16'h4E30: data_out = 8'h7E;
                    16'h4E31: data_out = 8'h7F;
                    16'h4E32: data_out = 8'h80;
                    16'h4E33: data_out = 8'h81;
                    16'h4E34: data_out = 8'h82;
                    16'h4E35: data_out = 8'h83;
                    16'h4E36: data_out = 8'h84;
                    16'h4E37: data_out = 8'h85;
                    16'h4E38: data_out = 8'h86;
                    16'h4E39: data_out = 8'h87;
                    16'h4E3A: data_out = 8'h88;
                    16'h4E3B: data_out = 8'h89;
                    16'h4E3C: data_out = 8'h8A;
                    16'h4E3D: data_out = 8'h8B;
                    16'h4E3E: data_out = 8'h8C;
                    16'h4E3F: data_out = 8'h8D;
                    16'h4E40: data_out = 8'h8E;
                    16'h4E41: data_out = 8'h8F;
                    16'h4E42: data_out = 8'h90;
                    16'h4E43: data_out = 8'h91;
                    16'h4E44: data_out = 8'h92;
                    16'h4E45: data_out = 8'h93;
                    16'h4E46: data_out = 8'h94;
                    16'h4E47: data_out = 8'h95;
                    16'h4E48: data_out = 8'h96;
                    16'h4E49: data_out = 8'h97;
                    16'h4E4A: data_out = 8'h98;
                    16'h4E4B: data_out = 8'h99;
                    16'h4E4C: data_out = 8'h9A;
                    16'h4E4D: data_out = 8'h9B;
                    16'h4E4E: data_out = 8'h9C;
                    16'h4E4F: data_out = 8'h9D;
                    16'h4E50: data_out = 8'h9E;
                    16'h4E51: data_out = 8'h9F;
                    16'h4E52: data_out = 8'hA0;
                    16'h4E53: data_out = 8'hA1;
                    16'h4E54: data_out = 8'hA2;
                    16'h4E55: data_out = 8'hA3;
                    16'h4E56: data_out = 8'hA4;
                    16'h4E57: data_out = 8'hA5;
                    16'h4E58: data_out = 8'hA6;
                    16'h4E59: data_out = 8'hA7;
                    16'h4E5A: data_out = 8'hA8;
                    16'h4E5B: data_out = 8'hA9;
                    16'h4E5C: data_out = 8'hAA;
                    16'h4E5D: data_out = 8'hAB;
                    16'h4E5E: data_out = 8'hAC;
                    16'h4E5F: data_out = 8'hAD;
                    16'h4E60: data_out = 8'hAE;
                    16'h4E61: data_out = 8'hAF;
                    16'h4E62: data_out = 8'hB0;
                    16'h4E63: data_out = 8'hB1;
                    16'h4E64: data_out = 8'hB2;
                    16'h4E65: data_out = 8'hB3;
                    16'h4E66: data_out = 8'hB4;
                    16'h4E67: data_out = 8'hB5;
                    16'h4E68: data_out = 8'hB6;
                    16'h4E69: data_out = 8'hB7;
                    16'h4E6A: data_out = 8'hB8;
                    16'h4E6B: data_out = 8'hB9;
                    16'h4E6C: data_out = 8'hBA;
                    16'h4E6D: data_out = 8'hBB;
                    16'h4E6E: data_out = 8'hBC;
                    16'h4E6F: data_out = 8'hBD;
                    16'h4E70: data_out = 8'hBE;
                    16'h4E71: data_out = 8'hBF;
                    16'h4E72: data_out = 8'hC0;
                    16'h4E73: data_out = 8'hC1;
                    16'h4E74: data_out = 8'hC2;
                    16'h4E75: data_out = 8'hC3;
                    16'h4E76: data_out = 8'hC4;
                    16'h4E77: data_out = 8'hC5;
                    16'h4E78: data_out = 8'hC6;
                    16'h4E79: data_out = 8'hC7;
                    16'h4E7A: data_out = 8'hC8;
                    16'h4E7B: data_out = 8'hC9;
                    16'h4E7C: data_out = 8'hCA;
                    16'h4E7D: data_out = 8'hCB;
                    16'h4E7E: data_out = 8'hCC;
                    16'h4E7F: data_out = 8'hCD;
                    16'h4E80: data_out = 8'h4E;
                    16'h4E81: data_out = 8'h4D;
                    16'h4E82: data_out = 8'h4C;
                    16'h4E83: data_out = 8'h4B;
                    16'h4E84: data_out = 8'h4A;
                    16'h4E85: data_out = 8'h49;
                    16'h4E86: data_out = 8'h48;
                    16'h4E87: data_out = 8'h47;
                    16'h4E88: data_out = 8'h46;
                    16'h4E89: data_out = 8'h45;
                    16'h4E8A: data_out = 8'h44;
                    16'h4E8B: data_out = 8'h43;
                    16'h4E8C: data_out = 8'h42;
                    16'h4E8D: data_out = 8'h41;
                    16'h4E8E: data_out = 8'h40;
                    16'h4E8F: data_out = 8'h3F;
                    16'h4E90: data_out = 8'h3E;
                    16'h4E91: data_out = 8'h3D;
                    16'h4E92: data_out = 8'h3C;
                    16'h4E93: data_out = 8'h3B;
                    16'h4E94: data_out = 8'h3A;
                    16'h4E95: data_out = 8'h39;
                    16'h4E96: data_out = 8'h38;
                    16'h4E97: data_out = 8'h37;
                    16'h4E98: data_out = 8'h36;
                    16'h4E99: data_out = 8'h35;
                    16'h4E9A: data_out = 8'h34;
                    16'h4E9B: data_out = 8'h33;
                    16'h4E9C: data_out = 8'h32;
                    16'h4E9D: data_out = 8'h31;
                    16'h4E9E: data_out = 8'h30;
                    16'h4E9F: data_out = 8'h2F;
                    16'h4EA0: data_out = 8'h2E;
                    16'h4EA1: data_out = 8'h2D;
                    16'h4EA2: data_out = 8'h2C;
                    16'h4EA3: data_out = 8'h2B;
                    16'h4EA4: data_out = 8'h2A;
                    16'h4EA5: data_out = 8'h29;
                    16'h4EA6: data_out = 8'h28;
                    16'h4EA7: data_out = 8'h27;
                    16'h4EA8: data_out = 8'h26;
                    16'h4EA9: data_out = 8'h25;
                    16'h4EAA: data_out = 8'h24;
                    16'h4EAB: data_out = 8'h23;
                    16'h4EAC: data_out = 8'h22;
                    16'h4EAD: data_out = 8'h21;
                    16'h4EAE: data_out = 8'h20;
                    16'h4EAF: data_out = 8'h1F;
                    16'h4EB0: data_out = 8'h1E;
                    16'h4EB1: data_out = 8'h1D;
                    16'h4EB2: data_out = 8'h1C;
                    16'h4EB3: data_out = 8'h1B;
                    16'h4EB4: data_out = 8'h1A;
                    16'h4EB5: data_out = 8'h19;
                    16'h4EB6: data_out = 8'h18;
                    16'h4EB7: data_out = 8'h17;
                    16'h4EB8: data_out = 8'h16;
                    16'h4EB9: data_out = 8'h15;
                    16'h4EBA: data_out = 8'h14;
                    16'h4EBB: data_out = 8'h13;
                    16'h4EBC: data_out = 8'h12;
                    16'h4EBD: data_out = 8'h11;
                    16'h4EBE: data_out = 8'h10;
                    16'h4EBF: data_out = 8'hF;
                    16'h4EC0: data_out = 8'hE;
                    16'h4EC1: data_out = 8'hD;
                    16'h4EC2: data_out = 8'hC;
                    16'h4EC3: data_out = 8'hB;
                    16'h4EC4: data_out = 8'hA;
                    16'h4EC5: data_out = 8'h9;
                    16'h4EC6: data_out = 8'h8;
                    16'h4EC7: data_out = 8'h7;
                    16'h4EC8: data_out = 8'h6;
                    16'h4EC9: data_out = 8'h5;
                    16'h4ECA: data_out = 8'h4;
                    16'h4ECB: data_out = 8'h3;
                    16'h4ECC: data_out = 8'h2;
                    16'h4ECD: data_out = 8'h1;
                    16'h4ECE: data_out = 8'h0;
                    16'h4ECF: data_out = 8'h81;
                    16'h4ED0: data_out = 8'h82;
                    16'h4ED1: data_out = 8'h83;
                    16'h4ED2: data_out = 8'h84;
                    16'h4ED3: data_out = 8'h85;
                    16'h4ED4: data_out = 8'h86;
                    16'h4ED5: data_out = 8'h87;
                    16'h4ED6: data_out = 8'h88;
                    16'h4ED7: data_out = 8'h89;
                    16'h4ED8: data_out = 8'h8A;
                    16'h4ED9: data_out = 8'h8B;
                    16'h4EDA: data_out = 8'h8C;
                    16'h4EDB: data_out = 8'h8D;
                    16'h4EDC: data_out = 8'h8E;
                    16'h4EDD: data_out = 8'h8F;
                    16'h4EDE: data_out = 8'h90;
                    16'h4EDF: data_out = 8'h91;
                    16'h4EE0: data_out = 8'h92;
                    16'h4EE1: data_out = 8'h93;
                    16'h4EE2: data_out = 8'h94;
                    16'h4EE3: data_out = 8'h95;
                    16'h4EE4: data_out = 8'h96;
                    16'h4EE5: data_out = 8'h97;
                    16'h4EE6: data_out = 8'h98;
                    16'h4EE7: data_out = 8'h99;
                    16'h4EE8: data_out = 8'h9A;
                    16'h4EE9: data_out = 8'h9B;
                    16'h4EEA: data_out = 8'h9C;
                    16'h4EEB: data_out = 8'h9D;
                    16'h4EEC: data_out = 8'h9E;
                    16'h4EED: data_out = 8'h9F;
                    16'h4EEE: data_out = 8'hA0;
                    16'h4EEF: data_out = 8'hA1;
                    16'h4EF0: data_out = 8'hA2;
                    16'h4EF1: data_out = 8'hA3;
                    16'h4EF2: data_out = 8'hA4;
                    16'h4EF3: data_out = 8'hA5;
                    16'h4EF4: data_out = 8'hA6;
                    16'h4EF5: data_out = 8'hA7;
                    16'h4EF6: data_out = 8'hA8;
                    16'h4EF7: data_out = 8'hA9;
                    16'h4EF8: data_out = 8'hAA;
                    16'h4EF9: data_out = 8'hAB;
                    16'h4EFA: data_out = 8'hAC;
                    16'h4EFB: data_out = 8'hAD;
                    16'h4EFC: data_out = 8'hAE;
                    16'h4EFD: data_out = 8'hAF;
                    16'h4EFE: data_out = 8'hB0;
                    16'h4EFF: data_out = 8'hB1;
                    16'h4F00: data_out = 8'h4F;
                    16'h4F01: data_out = 8'h50;
                    16'h4F02: data_out = 8'h51;
                    16'h4F03: data_out = 8'h52;
                    16'h4F04: data_out = 8'h53;
                    16'h4F05: data_out = 8'h54;
                    16'h4F06: data_out = 8'h55;
                    16'h4F07: data_out = 8'h56;
                    16'h4F08: data_out = 8'h57;
                    16'h4F09: data_out = 8'h58;
                    16'h4F0A: data_out = 8'h59;
                    16'h4F0B: data_out = 8'h5A;
                    16'h4F0C: data_out = 8'h5B;
                    16'h4F0D: data_out = 8'h5C;
                    16'h4F0E: data_out = 8'h5D;
                    16'h4F0F: data_out = 8'h5E;
                    16'h4F10: data_out = 8'h5F;
                    16'h4F11: data_out = 8'h60;
                    16'h4F12: data_out = 8'h61;
                    16'h4F13: data_out = 8'h62;
                    16'h4F14: data_out = 8'h63;
                    16'h4F15: data_out = 8'h64;
                    16'h4F16: data_out = 8'h65;
                    16'h4F17: data_out = 8'h66;
                    16'h4F18: data_out = 8'h67;
                    16'h4F19: data_out = 8'h68;
                    16'h4F1A: data_out = 8'h69;
                    16'h4F1B: data_out = 8'h6A;
                    16'h4F1C: data_out = 8'h6B;
                    16'h4F1D: data_out = 8'h6C;
                    16'h4F1E: data_out = 8'h6D;
                    16'h4F1F: data_out = 8'h6E;
                    16'h4F20: data_out = 8'h6F;
                    16'h4F21: data_out = 8'h70;
                    16'h4F22: data_out = 8'h71;
                    16'h4F23: data_out = 8'h72;
                    16'h4F24: data_out = 8'h73;
                    16'h4F25: data_out = 8'h74;
                    16'h4F26: data_out = 8'h75;
                    16'h4F27: data_out = 8'h76;
                    16'h4F28: data_out = 8'h77;
                    16'h4F29: data_out = 8'h78;
                    16'h4F2A: data_out = 8'h79;
                    16'h4F2B: data_out = 8'h7A;
                    16'h4F2C: data_out = 8'h7B;
                    16'h4F2D: data_out = 8'h7C;
                    16'h4F2E: data_out = 8'h7D;
                    16'h4F2F: data_out = 8'h7E;
                    16'h4F30: data_out = 8'h7F;
                    16'h4F31: data_out = 8'h80;
                    16'h4F32: data_out = 8'h81;
                    16'h4F33: data_out = 8'h82;
                    16'h4F34: data_out = 8'h83;
                    16'h4F35: data_out = 8'h84;
                    16'h4F36: data_out = 8'h85;
                    16'h4F37: data_out = 8'h86;
                    16'h4F38: data_out = 8'h87;
                    16'h4F39: data_out = 8'h88;
                    16'h4F3A: data_out = 8'h89;
                    16'h4F3B: data_out = 8'h8A;
                    16'h4F3C: data_out = 8'h8B;
                    16'h4F3D: data_out = 8'h8C;
                    16'h4F3E: data_out = 8'h8D;
                    16'h4F3F: data_out = 8'h8E;
                    16'h4F40: data_out = 8'h8F;
                    16'h4F41: data_out = 8'h90;
                    16'h4F42: data_out = 8'h91;
                    16'h4F43: data_out = 8'h92;
                    16'h4F44: data_out = 8'h93;
                    16'h4F45: data_out = 8'h94;
                    16'h4F46: data_out = 8'h95;
                    16'h4F47: data_out = 8'h96;
                    16'h4F48: data_out = 8'h97;
                    16'h4F49: data_out = 8'h98;
                    16'h4F4A: data_out = 8'h99;
                    16'h4F4B: data_out = 8'h9A;
                    16'h4F4C: data_out = 8'h9B;
                    16'h4F4D: data_out = 8'h9C;
                    16'h4F4E: data_out = 8'h9D;
                    16'h4F4F: data_out = 8'h9E;
                    16'h4F50: data_out = 8'h9F;
                    16'h4F51: data_out = 8'hA0;
                    16'h4F52: data_out = 8'hA1;
                    16'h4F53: data_out = 8'hA2;
                    16'h4F54: data_out = 8'hA3;
                    16'h4F55: data_out = 8'hA4;
                    16'h4F56: data_out = 8'hA5;
                    16'h4F57: data_out = 8'hA6;
                    16'h4F58: data_out = 8'hA7;
                    16'h4F59: data_out = 8'hA8;
                    16'h4F5A: data_out = 8'hA9;
                    16'h4F5B: data_out = 8'hAA;
                    16'h4F5C: data_out = 8'hAB;
                    16'h4F5D: data_out = 8'hAC;
                    16'h4F5E: data_out = 8'hAD;
                    16'h4F5F: data_out = 8'hAE;
                    16'h4F60: data_out = 8'hAF;
                    16'h4F61: data_out = 8'hB0;
                    16'h4F62: data_out = 8'hB1;
                    16'h4F63: data_out = 8'hB2;
                    16'h4F64: data_out = 8'hB3;
                    16'h4F65: data_out = 8'hB4;
                    16'h4F66: data_out = 8'hB5;
                    16'h4F67: data_out = 8'hB6;
                    16'h4F68: data_out = 8'hB7;
                    16'h4F69: data_out = 8'hB8;
                    16'h4F6A: data_out = 8'hB9;
                    16'h4F6B: data_out = 8'hBA;
                    16'h4F6C: data_out = 8'hBB;
                    16'h4F6D: data_out = 8'hBC;
                    16'h4F6E: data_out = 8'hBD;
                    16'h4F6F: data_out = 8'hBE;
                    16'h4F70: data_out = 8'hBF;
                    16'h4F71: data_out = 8'hC0;
                    16'h4F72: data_out = 8'hC1;
                    16'h4F73: data_out = 8'hC2;
                    16'h4F74: data_out = 8'hC3;
                    16'h4F75: data_out = 8'hC4;
                    16'h4F76: data_out = 8'hC5;
                    16'h4F77: data_out = 8'hC6;
                    16'h4F78: data_out = 8'hC7;
                    16'h4F79: data_out = 8'hC8;
                    16'h4F7A: data_out = 8'hC9;
                    16'h4F7B: data_out = 8'hCA;
                    16'h4F7C: data_out = 8'hCB;
                    16'h4F7D: data_out = 8'hCC;
                    16'h4F7E: data_out = 8'hCD;
                    16'h4F7F: data_out = 8'hCE;
                    16'h4F80: data_out = 8'h4F;
                    16'h4F81: data_out = 8'h4E;
                    16'h4F82: data_out = 8'h4D;
                    16'h4F83: data_out = 8'h4C;
                    16'h4F84: data_out = 8'h4B;
                    16'h4F85: data_out = 8'h4A;
                    16'h4F86: data_out = 8'h49;
                    16'h4F87: data_out = 8'h48;
                    16'h4F88: data_out = 8'h47;
                    16'h4F89: data_out = 8'h46;
                    16'h4F8A: data_out = 8'h45;
                    16'h4F8B: data_out = 8'h44;
                    16'h4F8C: data_out = 8'h43;
                    16'h4F8D: data_out = 8'h42;
                    16'h4F8E: data_out = 8'h41;
                    16'h4F8F: data_out = 8'h40;
                    16'h4F90: data_out = 8'h3F;
                    16'h4F91: data_out = 8'h3E;
                    16'h4F92: data_out = 8'h3D;
                    16'h4F93: data_out = 8'h3C;
                    16'h4F94: data_out = 8'h3B;
                    16'h4F95: data_out = 8'h3A;
                    16'h4F96: data_out = 8'h39;
                    16'h4F97: data_out = 8'h38;
                    16'h4F98: data_out = 8'h37;
                    16'h4F99: data_out = 8'h36;
                    16'h4F9A: data_out = 8'h35;
                    16'h4F9B: data_out = 8'h34;
                    16'h4F9C: data_out = 8'h33;
                    16'h4F9D: data_out = 8'h32;
                    16'h4F9E: data_out = 8'h31;
                    16'h4F9F: data_out = 8'h30;
                    16'h4FA0: data_out = 8'h2F;
                    16'h4FA1: data_out = 8'h2E;
                    16'h4FA2: data_out = 8'h2D;
                    16'h4FA3: data_out = 8'h2C;
                    16'h4FA4: data_out = 8'h2B;
                    16'h4FA5: data_out = 8'h2A;
                    16'h4FA6: data_out = 8'h29;
                    16'h4FA7: data_out = 8'h28;
                    16'h4FA8: data_out = 8'h27;
                    16'h4FA9: data_out = 8'h26;
                    16'h4FAA: data_out = 8'h25;
                    16'h4FAB: data_out = 8'h24;
                    16'h4FAC: data_out = 8'h23;
                    16'h4FAD: data_out = 8'h22;
                    16'h4FAE: data_out = 8'h21;
                    16'h4FAF: data_out = 8'h20;
                    16'h4FB0: data_out = 8'h1F;
                    16'h4FB1: data_out = 8'h1E;
                    16'h4FB2: data_out = 8'h1D;
                    16'h4FB3: data_out = 8'h1C;
                    16'h4FB4: data_out = 8'h1B;
                    16'h4FB5: data_out = 8'h1A;
                    16'h4FB6: data_out = 8'h19;
                    16'h4FB7: data_out = 8'h18;
                    16'h4FB8: data_out = 8'h17;
                    16'h4FB9: data_out = 8'h16;
                    16'h4FBA: data_out = 8'h15;
                    16'h4FBB: data_out = 8'h14;
                    16'h4FBC: data_out = 8'h13;
                    16'h4FBD: data_out = 8'h12;
                    16'h4FBE: data_out = 8'h11;
                    16'h4FBF: data_out = 8'h10;
                    16'h4FC0: data_out = 8'hF;
                    16'h4FC1: data_out = 8'hE;
                    16'h4FC2: data_out = 8'hD;
                    16'h4FC3: data_out = 8'hC;
                    16'h4FC4: data_out = 8'hB;
                    16'h4FC5: data_out = 8'hA;
                    16'h4FC6: data_out = 8'h9;
                    16'h4FC7: data_out = 8'h8;
                    16'h4FC8: data_out = 8'h7;
                    16'h4FC9: data_out = 8'h6;
                    16'h4FCA: data_out = 8'h5;
                    16'h4FCB: data_out = 8'h4;
                    16'h4FCC: data_out = 8'h3;
                    16'h4FCD: data_out = 8'h2;
                    16'h4FCE: data_out = 8'h1;
                    16'h4FCF: data_out = 8'h0;
                    16'h4FD0: data_out = 8'h81;
                    16'h4FD1: data_out = 8'h82;
                    16'h4FD2: data_out = 8'h83;
                    16'h4FD3: data_out = 8'h84;
                    16'h4FD4: data_out = 8'h85;
                    16'h4FD5: data_out = 8'h86;
                    16'h4FD6: data_out = 8'h87;
                    16'h4FD7: data_out = 8'h88;
                    16'h4FD8: data_out = 8'h89;
                    16'h4FD9: data_out = 8'h8A;
                    16'h4FDA: data_out = 8'h8B;
                    16'h4FDB: data_out = 8'h8C;
                    16'h4FDC: data_out = 8'h8D;
                    16'h4FDD: data_out = 8'h8E;
                    16'h4FDE: data_out = 8'h8F;
                    16'h4FDF: data_out = 8'h90;
                    16'h4FE0: data_out = 8'h91;
                    16'h4FE1: data_out = 8'h92;
                    16'h4FE2: data_out = 8'h93;
                    16'h4FE3: data_out = 8'h94;
                    16'h4FE4: data_out = 8'h95;
                    16'h4FE5: data_out = 8'h96;
                    16'h4FE6: data_out = 8'h97;
                    16'h4FE7: data_out = 8'h98;
                    16'h4FE8: data_out = 8'h99;
                    16'h4FE9: data_out = 8'h9A;
                    16'h4FEA: data_out = 8'h9B;
                    16'h4FEB: data_out = 8'h9C;
                    16'h4FEC: data_out = 8'h9D;
                    16'h4FED: data_out = 8'h9E;
                    16'h4FEE: data_out = 8'h9F;
                    16'h4FEF: data_out = 8'hA0;
                    16'h4FF0: data_out = 8'hA1;
                    16'h4FF1: data_out = 8'hA2;
                    16'h4FF2: data_out = 8'hA3;
                    16'h4FF3: data_out = 8'hA4;
                    16'h4FF4: data_out = 8'hA5;
                    16'h4FF5: data_out = 8'hA6;
                    16'h4FF6: data_out = 8'hA7;
                    16'h4FF7: data_out = 8'hA8;
                    16'h4FF8: data_out = 8'hA9;
                    16'h4FF9: data_out = 8'hAA;
                    16'h4FFA: data_out = 8'hAB;
                    16'h4FFB: data_out = 8'hAC;
                    16'h4FFC: data_out = 8'hAD;
                    16'h4FFD: data_out = 8'hAE;
                    16'h4FFE: data_out = 8'hAF;
                    16'h4FFF: data_out = 8'hB0;
                    16'h5000: data_out = 8'h50;
                    16'h5001: data_out = 8'h51;
                    16'h5002: data_out = 8'h52;
                    16'h5003: data_out = 8'h53;
                    16'h5004: data_out = 8'h54;
                    16'h5005: data_out = 8'h55;
                    16'h5006: data_out = 8'h56;
                    16'h5007: data_out = 8'h57;
                    16'h5008: data_out = 8'h58;
                    16'h5009: data_out = 8'h59;
                    16'h500A: data_out = 8'h5A;
                    16'h500B: data_out = 8'h5B;
                    16'h500C: data_out = 8'h5C;
                    16'h500D: data_out = 8'h5D;
                    16'h500E: data_out = 8'h5E;
                    16'h500F: data_out = 8'h5F;
                    16'h5010: data_out = 8'h60;
                    16'h5011: data_out = 8'h61;
                    16'h5012: data_out = 8'h62;
                    16'h5013: data_out = 8'h63;
                    16'h5014: data_out = 8'h64;
                    16'h5015: data_out = 8'h65;
                    16'h5016: data_out = 8'h66;
                    16'h5017: data_out = 8'h67;
                    16'h5018: data_out = 8'h68;
                    16'h5019: data_out = 8'h69;
                    16'h501A: data_out = 8'h6A;
                    16'h501B: data_out = 8'h6B;
                    16'h501C: data_out = 8'h6C;
                    16'h501D: data_out = 8'h6D;
                    16'h501E: data_out = 8'h6E;
                    16'h501F: data_out = 8'h6F;
                    16'h5020: data_out = 8'h70;
                    16'h5021: data_out = 8'h71;
                    16'h5022: data_out = 8'h72;
                    16'h5023: data_out = 8'h73;
                    16'h5024: data_out = 8'h74;
                    16'h5025: data_out = 8'h75;
                    16'h5026: data_out = 8'h76;
                    16'h5027: data_out = 8'h77;
                    16'h5028: data_out = 8'h78;
                    16'h5029: data_out = 8'h79;
                    16'h502A: data_out = 8'h7A;
                    16'h502B: data_out = 8'h7B;
                    16'h502C: data_out = 8'h7C;
                    16'h502D: data_out = 8'h7D;
                    16'h502E: data_out = 8'h7E;
                    16'h502F: data_out = 8'h7F;
                    16'h5030: data_out = 8'h80;
                    16'h5031: data_out = 8'h81;
                    16'h5032: data_out = 8'h82;
                    16'h5033: data_out = 8'h83;
                    16'h5034: data_out = 8'h84;
                    16'h5035: data_out = 8'h85;
                    16'h5036: data_out = 8'h86;
                    16'h5037: data_out = 8'h87;
                    16'h5038: data_out = 8'h88;
                    16'h5039: data_out = 8'h89;
                    16'h503A: data_out = 8'h8A;
                    16'h503B: data_out = 8'h8B;
                    16'h503C: data_out = 8'h8C;
                    16'h503D: data_out = 8'h8D;
                    16'h503E: data_out = 8'h8E;
                    16'h503F: data_out = 8'h8F;
                    16'h5040: data_out = 8'h90;
                    16'h5041: data_out = 8'h91;
                    16'h5042: data_out = 8'h92;
                    16'h5043: data_out = 8'h93;
                    16'h5044: data_out = 8'h94;
                    16'h5045: data_out = 8'h95;
                    16'h5046: data_out = 8'h96;
                    16'h5047: data_out = 8'h97;
                    16'h5048: data_out = 8'h98;
                    16'h5049: data_out = 8'h99;
                    16'h504A: data_out = 8'h9A;
                    16'h504B: data_out = 8'h9B;
                    16'h504C: data_out = 8'h9C;
                    16'h504D: data_out = 8'h9D;
                    16'h504E: data_out = 8'h9E;
                    16'h504F: data_out = 8'h9F;
                    16'h5050: data_out = 8'hA0;
                    16'h5051: data_out = 8'hA1;
                    16'h5052: data_out = 8'hA2;
                    16'h5053: data_out = 8'hA3;
                    16'h5054: data_out = 8'hA4;
                    16'h5055: data_out = 8'hA5;
                    16'h5056: data_out = 8'hA6;
                    16'h5057: data_out = 8'hA7;
                    16'h5058: data_out = 8'hA8;
                    16'h5059: data_out = 8'hA9;
                    16'h505A: data_out = 8'hAA;
                    16'h505B: data_out = 8'hAB;
                    16'h505C: data_out = 8'hAC;
                    16'h505D: data_out = 8'hAD;
                    16'h505E: data_out = 8'hAE;
                    16'h505F: data_out = 8'hAF;
                    16'h5060: data_out = 8'hB0;
                    16'h5061: data_out = 8'hB1;
                    16'h5062: data_out = 8'hB2;
                    16'h5063: data_out = 8'hB3;
                    16'h5064: data_out = 8'hB4;
                    16'h5065: data_out = 8'hB5;
                    16'h5066: data_out = 8'hB6;
                    16'h5067: data_out = 8'hB7;
                    16'h5068: data_out = 8'hB8;
                    16'h5069: data_out = 8'hB9;
                    16'h506A: data_out = 8'hBA;
                    16'h506B: data_out = 8'hBB;
                    16'h506C: data_out = 8'hBC;
                    16'h506D: data_out = 8'hBD;
                    16'h506E: data_out = 8'hBE;
                    16'h506F: data_out = 8'hBF;
                    16'h5070: data_out = 8'hC0;
                    16'h5071: data_out = 8'hC1;
                    16'h5072: data_out = 8'hC2;
                    16'h5073: data_out = 8'hC3;
                    16'h5074: data_out = 8'hC4;
                    16'h5075: data_out = 8'hC5;
                    16'h5076: data_out = 8'hC6;
                    16'h5077: data_out = 8'hC7;
                    16'h5078: data_out = 8'hC8;
                    16'h5079: data_out = 8'hC9;
                    16'h507A: data_out = 8'hCA;
                    16'h507B: data_out = 8'hCB;
                    16'h507C: data_out = 8'hCC;
                    16'h507D: data_out = 8'hCD;
                    16'h507E: data_out = 8'hCE;
                    16'h507F: data_out = 8'hCF;
                    16'h5080: data_out = 8'h50;
                    16'h5081: data_out = 8'h4F;
                    16'h5082: data_out = 8'h4E;
                    16'h5083: data_out = 8'h4D;
                    16'h5084: data_out = 8'h4C;
                    16'h5085: data_out = 8'h4B;
                    16'h5086: data_out = 8'h4A;
                    16'h5087: data_out = 8'h49;
                    16'h5088: data_out = 8'h48;
                    16'h5089: data_out = 8'h47;
                    16'h508A: data_out = 8'h46;
                    16'h508B: data_out = 8'h45;
                    16'h508C: data_out = 8'h44;
                    16'h508D: data_out = 8'h43;
                    16'h508E: data_out = 8'h42;
                    16'h508F: data_out = 8'h41;
                    16'h5090: data_out = 8'h40;
                    16'h5091: data_out = 8'h3F;
                    16'h5092: data_out = 8'h3E;
                    16'h5093: data_out = 8'h3D;
                    16'h5094: data_out = 8'h3C;
                    16'h5095: data_out = 8'h3B;
                    16'h5096: data_out = 8'h3A;
                    16'h5097: data_out = 8'h39;
                    16'h5098: data_out = 8'h38;
                    16'h5099: data_out = 8'h37;
                    16'h509A: data_out = 8'h36;
                    16'h509B: data_out = 8'h35;
                    16'h509C: data_out = 8'h34;
                    16'h509D: data_out = 8'h33;
                    16'h509E: data_out = 8'h32;
                    16'h509F: data_out = 8'h31;
                    16'h50A0: data_out = 8'h30;
                    16'h50A1: data_out = 8'h2F;
                    16'h50A2: data_out = 8'h2E;
                    16'h50A3: data_out = 8'h2D;
                    16'h50A4: data_out = 8'h2C;
                    16'h50A5: data_out = 8'h2B;
                    16'h50A6: data_out = 8'h2A;
                    16'h50A7: data_out = 8'h29;
                    16'h50A8: data_out = 8'h28;
                    16'h50A9: data_out = 8'h27;
                    16'h50AA: data_out = 8'h26;
                    16'h50AB: data_out = 8'h25;
                    16'h50AC: data_out = 8'h24;
                    16'h50AD: data_out = 8'h23;
                    16'h50AE: data_out = 8'h22;
                    16'h50AF: data_out = 8'h21;
                    16'h50B0: data_out = 8'h20;
                    16'h50B1: data_out = 8'h1F;
                    16'h50B2: data_out = 8'h1E;
                    16'h50B3: data_out = 8'h1D;
                    16'h50B4: data_out = 8'h1C;
                    16'h50B5: data_out = 8'h1B;
                    16'h50B6: data_out = 8'h1A;
                    16'h50B7: data_out = 8'h19;
                    16'h50B8: data_out = 8'h18;
                    16'h50B9: data_out = 8'h17;
                    16'h50BA: data_out = 8'h16;
                    16'h50BB: data_out = 8'h15;
                    16'h50BC: data_out = 8'h14;
                    16'h50BD: data_out = 8'h13;
                    16'h50BE: data_out = 8'h12;
                    16'h50BF: data_out = 8'h11;
                    16'h50C0: data_out = 8'h10;
                    16'h50C1: data_out = 8'hF;
                    16'h50C2: data_out = 8'hE;
                    16'h50C3: data_out = 8'hD;
                    16'h50C4: data_out = 8'hC;
                    16'h50C5: data_out = 8'hB;
                    16'h50C6: data_out = 8'hA;
                    16'h50C7: data_out = 8'h9;
                    16'h50C8: data_out = 8'h8;
                    16'h50C9: data_out = 8'h7;
                    16'h50CA: data_out = 8'h6;
                    16'h50CB: data_out = 8'h5;
                    16'h50CC: data_out = 8'h4;
                    16'h50CD: data_out = 8'h3;
                    16'h50CE: data_out = 8'h2;
                    16'h50CF: data_out = 8'h1;
                    16'h50D0: data_out = 8'h0;
                    16'h50D1: data_out = 8'h81;
                    16'h50D2: data_out = 8'h82;
                    16'h50D3: data_out = 8'h83;
                    16'h50D4: data_out = 8'h84;
                    16'h50D5: data_out = 8'h85;
                    16'h50D6: data_out = 8'h86;
                    16'h50D7: data_out = 8'h87;
                    16'h50D8: data_out = 8'h88;
                    16'h50D9: data_out = 8'h89;
                    16'h50DA: data_out = 8'h8A;
                    16'h50DB: data_out = 8'h8B;
                    16'h50DC: data_out = 8'h8C;
                    16'h50DD: data_out = 8'h8D;
                    16'h50DE: data_out = 8'h8E;
                    16'h50DF: data_out = 8'h8F;
                    16'h50E0: data_out = 8'h90;
                    16'h50E1: data_out = 8'h91;
                    16'h50E2: data_out = 8'h92;
                    16'h50E3: data_out = 8'h93;
                    16'h50E4: data_out = 8'h94;
                    16'h50E5: data_out = 8'h95;
                    16'h50E6: data_out = 8'h96;
                    16'h50E7: data_out = 8'h97;
                    16'h50E8: data_out = 8'h98;
                    16'h50E9: data_out = 8'h99;
                    16'h50EA: data_out = 8'h9A;
                    16'h50EB: data_out = 8'h9B;
                    16'h50EC: data_out = 8'h9C;
                    16'h50ED: data_out = 8'h9D;
                    16'h50EE: data_out = 8'h9E;
                    16'h50EF: data_out = 8'h9F;
                    16'h50F0: data_out = 8'hA0;
                    16'h50F1: data_out = 8'hA1;
                    16'h50F2: data_out = 8'hA2;
                    16'h50F3: data_out = 8'hA3;
                    16'h50F4: data_out = 8'hA4;
                    16'h50F5: data_out = 8'hA5;
                    16'h50F6: data_out = 8'hA6;
                    16'h50F7: data_out = 8'hA7;
                    16'h50F8: data_out = 8'hA8;
                    16'h50F9: data_out = 8'hA9;
                    16'h50FA: data_out = 8'hAA;
                    16'h50FB: data_out = 8'hAB;
                    16'h50FC: data_out = 8'hAC;
                    16'h50FD: data_out = 8'hAD;
                    16'h50FE: data_out = 8'hAE;
                    16'h50FF: data_out = 8'hAF;
                    16'h5100: data_out = 8'h51;
                    16'h5101: data_out = 8'h52;
                    16'h5102: data_out = 8'h53;
                    16'h5103: data_out = 8'h54;
                    16'h5104: data_out = 8'h55;
                    16'h5105: data_out = 8'h56;
                    16'h5106: data_out = 8'h57;
                    16'h5107: data_out = 8'h58;
                    16'h5108: data_out = 8'h59;
                    16'h5109: data_out = 8'h5A;
                    16'h510A: data_out = 8'h5B;
                    16'h510B: data_out = 8'h5C;
                    16'h510C: data_out = 8'h5D;
                    16'h510D: data_out = 8'h5E;
                    16'h510E: data_out = 8'h5F;
                    16'h510F: data_out = 8'h60;
                    16'h5110: data_out = 8'h61;
                    16'h5111: data_out = 8'h62;
                    16'h5112: data_out = 8'h63;
                    16'h5113: data_out = 8'h64;
                    16'h5114: data_out = 8'h65;
                    16'h5115: data_out = 8'h66;
                    16'h5116: data_out = 8'h67;
                    16'h5117: data_out = 8'h68;
                    16'h5118: data_out = 8'h69;
                    16'h5119: data_out = 8'h6A;
                    16'h511A: data_out = 8'h6B;
                    16'h511B: data_out = 8'h6C;
                    16'h511C: data_out = 8'h6D;
                    16'h511D: data_out = 8'h6E;
                    16'h511E: data_out = 8'h6F;
                    16'h511F: data_out = 8'h70;
                    16'h5120: data_out = 8'h71;
                    16'h5121: data_out = 8'h72;
                    16'h5122: data_out = 8'h73;
                    16'h5123: data_out = 8'h74;
                    16'h5124: data_out = 8'h75;
                    16'h5125: data_out = 8'h76;
                    16'h5126: data_out = 8'h77;
                    16'h5127: data_out = 8'h78;
                    16'h5128: data_out = 8'h79;
                    16'h5129: data_out = 8'h7A;
                    16'h512A: data_out = 8'h7B;
                    16'h512B: data_out = 8'h7C;
                    16'h512C: data_out = 8'h7D;
                    16'h512D: data_out = 8'h7E;
                    16'h512E: data_out = 8'h7F;
                    16'h512F: data_out = 8'h80;
                    16'h5130: data_out = 8'h81;
                    16'h5131: data_out = 8'h82;
                    16'h5132: data_out = 8'h83;
                    16'h5133: data_out = 8'h84;
                    16'h5134: data_out = 8'h85;
                    16'h5135: data_out = 8'h86;
                    16'h5136: data_out = 8'h87;
                    16'h5137: data_out = 8'h88;
                    16'h5138: data_out = 8'h89;
                    16'h5139: data_out = 8'h8A;
                    16'h513A: data_out = 8'h8B;
                    16'h513B: data_out = 8'h8C;
                    16'h513C: data_out = 8'h8D;
                    16'h513D: data_out = 8'h8E;
                    16'h513E: data_out = 8'h8F;
                    16'h513F: data_out = 8'h90;
                    16'h5140: data_out = 8'h91;
                    16'h5141: data_out = 8'h92;
                    16'h5142: data_out = 8'h93;
                    16'h5143: data_out = 8'h94;
                    16'h5144: data_out = 8'h95;
                    16'h5145: data_out = 8'h96;
                    16'h5146: data_out = 8'h97;
                    16'h5147: data_out = 8'h98;
                    16'h5148: data_out = 8'h99;
                    16'h5149: data_out = 8'h9A;
                    16'h514A: data_out = 8'h9B;
                    16'h514B: data_out = 8'h9C;
                    16'h514C: data_out = 8'h9D;
                    16'h514D: data_out = 8'h9E;
                    16'h514E: data_out = 8'h9F;
                    16'h514F: data_out = 8'hA0;
                    16'h5150: data_out = 8'hA1;
                    16'h5151: data_out = 8'hA2;
                    16'h5152: data_out = 8'hA3;
                    16'h5153: data_out = 8'hA4;
                    16'h5154: data_out = 8'hA5;
                    16'h5155: data_out = 8'hA6;
                    16'h5156: data_out = 8'hA7;
                    16'h5157: data_out = 8'hA8;
                    16'h5158: data_out = 8'hA9;
                    16'h5159: data_out = 8'hAA;
                    16'h515A: data_out = 8'hAB;
                    16'h515B: data_out = 8'hAC;
                    16'h515C: data_out = 8'hAD;
                    16'h515D: data_out = 8'hAE;
                    16'h515E: data_out = 8'hAF;
                    16'h515F: data_out = 8'hB0;
                    16'h5160: data_out = 8'hB1;
                    16'h5161: data_out = 8'hB2;
                    16'h5162: data_out = 8'hB3;
                    16'h5163: data_out = 8'hB4;
                    16'h5164: data_out = 8'hB5;
                    16'h5165: data_out = 8'hB6;
                    16'h5166: data_out = 8'hB7;
                    16'h5167: data_out = 8'hB8;
                    16'h5168: data_out = 8'hB9;
                    16'h5169: data_out = 8'hBA;
                    16'h516A: data_out = 8'hBB;
                    16'h516B: data_out = 8'hBC;
                    16'h516C: data_out = 8'hBD;
                    16'h516D: data_out = 8'hBE;
                    16'h516E: data_out = 8'hBF;
                    16'h516F: data_out = 8'hC0;
                    16'h5170: data_out = 8'hC1;
                    16'h5171: data_out = 8'hC2;
                    16'h5172: data_out = 8'hC3;
                    16'h5173: data_out = 8'hC4;
                    16'h5174: data_out = 8'hC5;
                    16'h5175: data_out = 8'hC6;
                    16'h5176: data_out = 8'hC7;
                    16'h5177: data_out = 8'hC8;
                    16'h5178: data_out = 8'hC9;
                    16'h5179: data_out = 8'hCA;
                    16'h517A: data_out = 8'hCB;
                    16'h517B: data_out = 8'hCC;
                    16'h517C: data_out = 8'hCD;
                    16'h517D: data_out = 8'hCE;
                    16'h517E: data_out = 8'hCF;
                    16'h517F: data_out = 8'hD0;
                    16'h5180: data_out = 8'h51;
                    16'h5181: data_out = 8'h50;
                    16'h5182: data_out = 8'h4F;
                    16'h5183: data_out = 8'h4E;
                    16'h5184: data_out = 8'h4D;
                    16'h5185: data_out = 8'h4C;
                    16'h5186: data_out = 8'h4B;
                    16'h5187: data_out = 8'h4A;
                    16'h5188: data_out = 8'h49;
                    16'h5189: data_out = 8'h48;
                    16'h518A: data_out = 8'h47;
                    16'h518B: data_out = 8'h46;
                    16'h518C: data_out = 8'h45;
                    16'h518D: data_out = 8'h44;
                    16'h518E: data_out = 8'h43;
                    16'h518F: data_out = 8'h42;
                    16'h5190: data_out = 8'h41;
                    16'h5191: data_out = 8'h40;
                    16'h5192: data_out = 8'h3F;
                    16'h5193: data_out = 8'h3E;
                    16'h5194: data_out = 8'h3D;
                    16'h5195: data_out = 8'h3C;
                    16'h5196: data_out = 8'h3B;
                    16'h5197: data_out = 8'h3A;
                    16'h5198: data_out = 8'h39;
                    16'h5199: data_out = 8'h38;
                    16'h519A: data_out = 8'h37;
                    16'h519B: data_out = 8'h36;
                    16'h519C: data_out = 8'h35;
                    16'h519D: data_out = 8'h34;
                    16'h519E: data_out = 8'h33;
                    16'h519F: data_out = 8'h32;
                    16'h51A0: data_out = 8'h31;
                    16'h51A1: data_out = 8'h30;
                    16'h51A2: data_out = 8'h2F;
                    16'h51A3: data_out = 8'h2E;
                    16'h51A4: data_out = 8'h2D;
                    16'h51A5: data_out = 8'h2C;
                    16'h51A6: data_out = 8'h2B;
                    16'h51A7: data_out = 8'h2A;
                    16'h51A8: data_out = 8'h29;
                    16'h51A9: data_out = 8'h28;
                    16'h51AA: data_out = 8'h27;
                    16'h51AB: data_out = 8'h26;
                    16'h51AC: data_out = 8'h25;
                    16'h51AD: data_out = 8'h24;
                    16'h51AE: data_out = 8'h23;
                    16'h51AF: data_out = 8'h22;
                    16'h51B0: data_out = 8'h21;
                    16'h51B1: data_out = 8'h20;
                    16'h51B2: data_out = 8'h1F;
                    16'h51B3: data_out = 8'h1E;
                    16'h51B4: data_out = 8'h1D;
                    16'h51B5: data_out = 8'h1C;
                    16'h51B6: data_out = 8'h1B;
                    16'h51B7: data_out = 8'h1A;
                    16'h51B8: data_out = 8'h19;
                    16'h51B9: data_out = 8'h18;
                    16'h51BA: data_out = 8'h17;
                    16'h51BB: data_out = 8'h16;
                    16'h51BC: data_out = 8'h15;
                    16'h51BD: data_out = 8'h14;
                    16'h51BE: data_out = 8'h13;
                    16'h51BF: data_out = 8'h12;
                    16'h51C0: data_out = 8'h11;
                    16'h51C1: data_out = 8'h10;
                    16'h51C2: data_out = 8'hF;
                    16'h51C3: data_out = 8'hE;
                    16'h51C4: data_out = 8'hD;
                    16'h51C5: data_out = 8'hC;
                    16'h51C6: data_out = 8'hB;
                    16'h51C7: data_out = 8'hA;
                    16'h51C8: data_out = 8'h9;
                    16'h51C9: data_out = 8'h8;
                    16'h51CA: data_out = 8'h7;
                    16'h51CB: data_out = 8'h6;
                    16'h51CC: data_out = 8'h5;
                    16'h51CD: data_out = 8'h4;
                    16'h51CE: data_out = 8'h3;
                    16'h51CF: data_out = 8'h2;
                    16'h51D0: data_out = 8'h1;
                    16'h51D1: data_out = 8'h0;
                    16'h51D2: data_out = 8'h81;
                    16'h51D3: data_out = 8'h82;
                    16'h51D4: data_out = 8'h83;
                    16'h51D5: data_out = 8'h84;
                    16'h51D6: data_out = 8'h85;
                    16'h51D7: data_out = 8'h86;
                    16'h51D8: data_out = 8'h87;
                    16'h51D9: data_out = 8'h88;
                    16'h51DA: data_out = 8'h89;
                    16'h51DB: data_out = 8'h8A;
                    16'h51DC: data_out = 8'h8B;
                    16'h51DD: data_out = 8'h8C;
                    16'h51DE: data_out = 8'h8D;
                    16'h51DF: data_out = 8'h8E;
                    16'h51E0: data_out = 8'h8F;
                    16'h51E1: data_out = 8'h90;
                    16'h51E2: data_out = 8'h91;
                    16'h51E3: data_out = 8'h92;
                    16'h51E4: data_out = 8'h93;
                    16'h51E5: data_out = 8'h94;
                    16'h51E6: data_out = 8'h95;
                    16'h51E7: data_out = 8'h96;
                    16'h51E8: data_out = 8'h97;
                    16'h51E9: data_out = 8'h98;
                    16'h51EA: data_out = 8'h99;
                    16'h51EB: data_out = 8'h9A;
                    16'h51EC: data_out = 8'h9B;
                    16'h51ED: data_out = 8'h9C;
                    16'h51EE: data_out = 8'h9D;
                    16'h51EF: data_out = 8'h9E;
                    16'h51F0: data_out = 8'h9F;
                    16'h51F1: data_out = 8'hA0;
                    16'h51F2: data_out = 8'hA1;
                    16'h51F3: data_out = 8'hA2;
                    16'h51F4: data_out = 8'hA3;
                    16'h51F5: data_out = 8'hA4;
                    16'h51F6: data_out = 8'hA5;
                    16'h51F7: data_out = 8'hA6;
                    16'h51F8: data_out = 8'hA7;
                    16'h51F9: data_out = 8'hA8;
                    16'h51FA: data_out = 8'hA9;
                    16'h51FB: data_out = 8'hAA;
                    16'h51FC: data_out = 8'hAB;
                    16'h51FD: data_out = 8'hAC;
                    16'h51FE: data_out = 8'hAD;
                    16'h51FF: data_out = 8'hAE;
                    16'h5200: data_out = 8'h52;
                    16'h5201: data_out = 8'h53;
                    16'h5202: data_out = 8'h54;
                    16'h5203: data_out = 8'h55;
                    16'h5204: data_out = 8'h56;
                    16'h5205: data_out = 8'h57;
                    16'h5206: data_out = 8'h58;
                    16'h5207: data_out = 8'h59;
                    16'h5208: data_out = 8'h5A;
                    16'h5209: data_out = 8'h5B;
                    16'h520A: data_out = 8'h5C;
                    16'h520B: data_out = 8'h5D;
                    16'h520C: data_out = 8'h5E;
                    16'h520D: data_out = 8'h5F;
                    16'h520E: data_out = 8'h60;
                    16'h520F: data_out = 8'h61;
                    16'h5210: data_out = 8'h62;
                    16'h5211: data_out = 8'h63;
                    16'h5212: data_out = 8'h64;
                    16'h5213: data_out = 8'h65;
                    16'h5214: data_out = 8'h66;
                    16'h5215: data_out = 8'h67;
                    16'h5216: data_out = 8'h68;
                    16'h5217: data_out = 8'h69;
                    16'h5218: data_out = 8'h6A;
                    16'h5219: data_out = 8'h6B;
                    16'h521A: data_out = 8'h6C;
                    16'h521B: data_out = 8'h6D;
                    16'h521C: data_out = 8'h6E;
                    16'h521D: data_out = 8'h6F;
                    16'h521E: data_out = 8'h70;
                    16'h521F: data_out = 8'h71;
                    16'h5220: data_out = 8'h72;
                    16'h5221: data_out = 8'h73;
                    16'h5222: data_out = 8'h74;
                    16'h5223: data_out = 8'h75;
                    16'h5224: data_out = 8'h76;
                    16'h5225: data_out = 8'h77;
                    16'h5226: data_out = 8'h78;
                    16'h5227: data_out = 8'h79;
                    16'h5228: data_out = 8'h7A;
                    16'h5229: data_out = 8'h7B;
                    16'h522A: data_out = 8'h7C;
                    16'h522B: data_out = 8'h7D;
                    16'h522C: data_out = 8'h7E;
                    16'h522D: data_out = 8'h7F;
                    16'h522E: data_out = 8'h80;
                    16'h522F: data_out = 8'h81;
                    16'h5230: data_out = 8'h82;
                    16'h5231: data_out = 8'h83;
                    16'h5232: data_out = 8'h84;
                    16'h5233: data_out = 8'h85;
                    16'h5234: data_out = 8'h86;
                    16'h5235: data_out = 8'h87;
                    16'h5236: data_out = 8'h88;
                    16'h5237: data_out = 8'h89;
                    16'h5238: data_out = 8'h8A;
                    16'h5239: data_out = 8'h8B;
                    16'h523A: data_out = 8'h8C;
                    16'h523B: data_out = 8'h8D;
                    16'h523C: data_out = 8'h8E;
                    16'h523D: data_out = 8'h8F;
                    16'h523E: data_out = 8'h90;
                    16'h523F: data_out = 8'h91;
                    16'h5240: data_out = 8'h92;
                    16'h5241: data_out = 8'h93;
                    16'h5242: data_out = 8'h94;
                    16'h5243: data_out = 8'h95;
                    16'h5244: data_out = 8'h96;
                    16'h5245: data_out = 8'h97;
                    16'h5246: data_out = 8'h98;
                    16'h5247: data_out = 8'h99;
                    16'h5248: data_out = 8'h9A;
                    16'h5249: data_out = 8'h9B;
                    16'h524A: data_out = 8'h9C;
                    16'h524B: data_out = 8'h9D;
                    16'h524C: data_out = 8'h9E;
                    16'h524D: data_out = 8'h9F;
                    16'h524E: data_out = 8'hA0;
                    16'h524F: data_out = 8'hA1;
                    16'h5250: data_out = 8'hA2;
                    16'h5251: data_out = 8'hA3;
                    16'h5252: data_out = 8'hA4;
                    16'h5253: data_out = 8'hA5;
                    16'h5254: data_out = 8'hA6;
                    16'h5255: data_out = 8'hA7;
                    16'h5256: data_out = 8'hA8;
                    16'h5257: data_out = 8'hA9;
                    16'h5258: data_out = 8'hAA;
                    16'h5259: data_out = 8'hAB;
                    16'h525A: data_out = 8'hAC;
                    16'h525B: data_out = 8'hAD;
                    16'h525C: data_out = 8'hAE;
                    16'h525D: data_out = 8'hAF;
                    16'h525E: data_out = 8'hB0;
                    16'h525F: data_out = 8'hB1;
                    16'h5260: data_out = 8'hB2;
                    16'h5261: data_out = 8'hB3;
                    16'h5262: data_out = 8'hB4;
                    16'h5263: data_out = 8'hB5;
                    16'h5264: data_out = 8'hB6;
                    16'h5265: data_out = 8'hB7;
                    16'h5266: data_out = 8'hB8;
                    16'h5267: data_out = 8'hB9;
                    16'h5268: data_out = 8'hBA;
                    16'h5269: data_out = 8'hBB;
                    16'h526A: data_out = 8'hBC;
                    16'h526B: data_out = 8'hBD;
                    16'h526C: data_out = 8'hBE;
                    16'h526D: data_out = 8'hBF;
                    16'h526E: data_out = 8'hC0;
                    16'h526F: data_out = 8'hC1;
                    16'h5270: data_out = 8'hC2;
                    16'h5271: data_out = 8'hC3;
                    16'h5272: data_out = 8'hC4;
                    16'h5273: data_out = 8'hC5;
                    16'h5274: data_out = 8'hC6;
                    16'h5275: data_out = 8'hC7;
                    16'h5276: data_out = 8'hC8;
                    16'h5277: data_out = 8'hC9;
                    16'h5278: data_out = 8'hCA;
                    16'h5279: data_out = 8'hCB;
                    16'h527A: data_out = 8'hCC;
                    16'h527B: data_out = 8'hCD;
                    16'h527C: data_out = 8'hCE;
                    16'h527D: data_out = 8'hCF;
                    16'h527E: data_out = 8'hD0;
                    16'h527F: data_out = 8'hD1;
                    16'h5280: data_out = 8'h52;
                    16'h5281: data_out = 8'h51;
                    16'h5282: data_out = 8'h50;
                    16'h5283: data_out = 8'h4F;
                    16'h5284: data_out = 8'h4E;
                    16'h5285: data_out = 8'h4D;
                    16'h5286: data_out = 8'h4C;
                    16'h5287: data_out = 8'h4B;
                    16'h5288: data_out = 8'h4A;
                    16'h5289: data_out = 8'h49;
                    16'h528A: data_out = 8'h48;
                    16'h528B: data_out = 8'h47;
                    16'h528C: data_out = 8'h46;
                    16'h528D: data_out = 8'h45;
                    16'h528E: data_out = 8'h44;
                    16'h528F: data_out = 8'h43;
                    16'h5290: data_out = 8'h42;
                    16'h5291: data_out = 8'h41;
                    16'h5292: data_out = 8'h40;
                    16'h5293: data_out = 8'h3F;
                    16'h5294: data_out = 8'h3E;
                    16'h5295: data_out = 8'h3D;
                    16'h5296: data_out = 8'h3C;
                    16'h5297: data_out = 8'h3B;
                    16'h5298: data_out = 8'h3A;
                    16'h5299: data_out = 8'h39;
                    16'h529A: data_out = 8'h38;
                    16'h529B: data_out = 8'h37;
                    16'h529C: data_out = 8'h36;
                    16'h529D: data_out = 8'h35;
                    16'h529E: data_out = 8'h34;
                    16'h529F: data_out = 8'h33;
                    16'h52A0: data_out = 8'h32;
                    16'h52A1: data_out = 8'h31;
                    16'h52A2: data_out = 8'h30;
                    16'h52A3: data_out = 8'h2F;
                    16'h52A4: data_out = 8'h2E;
                    16'h52A5: data_out = 8'h2D;
                    16'h52A6: data_out = 8'h2C;
                    16'h52A7: data_out = 8'h2B;
                    16'h52A8: data_out = 8'h2A;
                    16'h52A9: data_out = 8'h29;
                    16'h52AA: data_out = 8'h28;
                    16'h52AB: data_out = 8'h27;
                    16'h52AC: data_out = 8'h26;
                    16'h52AD: data_out = 8'h25;
                    16'h52AE: data_out = 8'h24;
                    16'h52AF: data_out = 8'h23;
                    16'h52B0: data_out = 8'h22;
                    16'h52B1: data_out = 8'h21;
                    16'h52B2: data_out = 8'h20;
                    16'h52B3: data_out = 8'h1F;
                    16'h52B4: data_out = 8'h1E;
                    16'h52B5: data_out = 8'h1D;
                    16'h52B6: data_out = 8'h1C;
                    16'h52B7: data_out = 8'h1B;
                    16'h52B8: data_out = 8'h1A;
                    16'h52B9: data_out = 8'h19;
                    16'h52BA: data_out = 8'h18;
                    16'h52BB: data_out = 8'h17;
                    16'h52BC: data_out = 8'h16;
                    16'h52BD: data_out = 8'h15;
                    16'h52BE: data_out = 8'h14;
                    16'h52BF: data_out = 8'h13;
                    16'h52C0: data_out = 8'h12;
                    16'h52C1: data_out = 8'h11;
                    16'h52C2: data_out = 8'h10;
                    16'h52C3: data_out = 8'hF;
                    16'h52C4: data_out = 8'hE;
                    16'h52C5: data_out = 8'hD;
                    16'h52C6: data_out = 8'hC;
                    16'h52C7: data_out = 8'hB;
                    16'h52C8: data_out = 8'hA;
                    16'h52C9: data_out = 8'h9;
                    16'h52CA: data_out = 8'h8;
                    16'h52CB: data_out = 8'h7;
                    16'h52CC: data_out = 8'h6;
                    16'h52CD: data_out = 8'h5;
                    16'h52CE: data_out = 8'h4;
                    16'h52CF: data_out = 8'h3;
                    16'h52D0: data_out = 8'h2;
                    16'h52D1: data_out = 8'h1;
                    16'h52D2: data_out = 8'h0;
                    16'h52D3: data_out = 8'h81;
                    16'h52D4: data_out = 8'h82;
                    16'h52D5: data_out = 8'h83;
                    16'h52D6: data_out = 8'h84;
                    16'h52D7: data_out = 8'h85;
                    16'h52D8: data_out = 8'h86;
                    16'h52D9: data_out = 8'h87;
                    16'h52DA: data_out = 8'h88;
                    16'h52DB: data_out = 8'h89;
                    16'h52DC: data_out = 8'h8A;
                    16'h52DD: data_out = 8'h8B;
                    16'h52DE: data_out = 8'h8C;
                    16'h52DF: data_out = 8'h8D;
                    16'h52E0: data_out = 8'h8E;
                    16'h52E1: data_out = 8'h8F;
                    16'h52E2: data_out = 8'h90;
                    16'h52E3: data_out = 8'h91;
                    16'h52E4: data_out = 8'h92;
                    16'h52E5: data_out = 8'h93;
                    16'h52E6: data_out = 8'h94;
                    16'h52E7: data_out = 8'h95;
                    16'h52E8: data_out = 8'h96;
                    16'h52E9: data_out = 8'h97;
                    16'h52EA: data_out = 8'h98;
                    16'h52EB: data_out = 8'h99;
                    16'h52EC: data_out = 8'h9A;
                    16'h52ED: data_out = 8'h9B;
                    16'h52EE: data_out = 8'h9C;
                    16'h52EF: data_out = 8'h9D;
                    16'h52F0: data_out = 8'h9E;
                    16'h52F1: data_out = 8'h9F;
                    16'h52F2: data_out = 8'hA0;
                    16'h52F3: data_out = 8'hA1;
                    16'h52F4: data_out = 8'hA2;
                    16'h52F5: data_out = 8'hA3;
                    16'h52F6: data_out = 8'hA4;
                    16'h52F7: data_out = 8'hA5;
                    16'h52F8: data_out = 8'hA6;
                    16'h52F9: data_out = 8'hA7;
                    16'h52FA: data_out = 8'hA8;
                    16'h52FB: data_out = 8'hA9;
                    16'h52FC: data_out = 8'hAA;
                    16'h52FD: data_out = 8'hAB;
                    16'h52FE: data_out = 8'hAC;
                    16'h52FF: data_out = 8'hAD;
                    16'h5300: data_out = 8'h53;
                    16'h5301: data_out = 8'h54;
                    16'h5302: data_out = 8'h55;
                    16'h5303: data_out = 8'h56;
                    16'h5304: data_out = 8'h57;
                    16'h5305: data_out = 8'h58;
                    16'h5306: data_out = 8'h59;
                    16'h5307: data_out = 8'h5A;
                    16'h5308: data_out = 8'h5B;
                    16'h5309: data_out = 8'h5C;
                    16'h530A: data_out = 8'h5D;
                    16'h530B: data_out = 8'h5E;
                    16'h530C: data_out = 8'h5F;
                    16'h530D: data_out = 8'h60;
                    16'h530E: data_out = 8'h61;
                    16'h530F: data_out = 8'h62;
                    16'h5310: data_out = 8'h63;
                    16'h5311: data_out = 8'h64;
                    16'h5312: data_out = 8'h65;
                    16'h5313: data_out = 8'h66;
                    16'h5314: data_out = 8'h67;
                    16'h5315: data_out = 8'h68;
                    16'h5316: data_out = 8'h69;
                    16'h5317: data_out = 8'h6A;
                    16'h5318: data_out = 8'h6B;
                    16'h5319: data_out = 8'h6C;
                    16'h531A: data_out = 8'h6D;
                    16'h531B: data_out = 8'h6E;
                    16'h531C: data_out = 8'h6F;
                    16'h531D: data_out = 8'h70;
                    16'h531E: data_out = 8'h71;
                    16'h531F: data_out = 8'h72;
                    16'h5320: data_out = 8'h73;
                    16'h5321: data_out = 8'h74;
                    16'h5322: data_out = 8'h75;
                    16'h5323: data_out = 8'h76;
                    16'h5324: data_out = 8'h77;
                    16'h5325: data_out = 8'h78;
                    16'h5326: data_out = 8'h79;
                    16'h5327: data_out = 8'h7A;
                    16'h5328: data_out = 8'h7B;
                    16'h5329: data_out = 8'h7C;
                    16'h532A: data_out = 8'h7D;
                    16'h532B: data_out = 8'h7E;
                    16'h532C: data_out = 8'h7F;
                    16'h532D: data_out = 8'h80;
                    16'h532E: data_out = 8'h81;
                    16'h532F: data_out = 8'h82;
                    16'h5330: data_out = 8'h83;
                    16'h5331: data_out = 8'h84;
                    16'h5332: data_out = 8'h85;
                    16'h5333: data_out = 8'h86;
                    16'h5334: data_out = 8'h87;
                    16'h5335: data_out = 8'h88;
                    16'h5336: data_out = 8'h89;
                    16'h5337: data_out = 8'h8A;
                    16'h5338: data_out = 8'h8B;
                    16'h5339: data_out = 8'h8C;
                    16'h533A: data_out = 8'h8D;
                    16'h533B: data_out = 8'h8E;
                    16'h533C: data_out = 8'h8F;
                    16'h533D: data_out = 8'h90;
                    16'h533E: data_out = 8'h91;
                    16'h533F: data_out = 8'h92;
                    16'h5340: data_out = 8'h93;
                    16'h5341: data_out = 8'h94;
                    16'h5342: data_out = 8'h95;
                    16'h5343: data_out = 8'h96;
                    16'h5344: data_out = 8'h97;
                    16'h5345: data_out = 8'h98;
                    16'h5346: data_out = 8'h99;
                    16'h5347: data_out = 8'h9A;
                    16'h5348: data_out = 8'h9B;
                    16'h5349: data_out = 8'h9C;
                    16'h534A: data_out = 8'h9D;
                    16'h534B: data_out = 8'h9E;
                    16'h534C: data_out = 8'h9F;
                    16'h534D: data_out = 8'hA0;
                    16'h534E: data_out = 8'hA1;
                    16'h534F: data_out = 8'hA2;
                    16'h5350: data_out = 8'hA3;
                    16'h5351: data_out = 8'hA4;
                    16'h5352: data_out = 8'hA5;
                    16'h5353: data_out = 8'hA6;
                    16'h5354: data_out = 8'hA7;
                    16'h5355: data_out = 8'hA8;
                    16'h5356: data_out = 8'hA9;
                    16'h5357: data_out = 8'hAA;
                    16'h5358: data_out = 8'hAB;
                    16'h5359: data_out = 8'hAC;
                    16'h535A: data_out = 8'hAD;
                    16'h535B: data_out = 8'hAE;
                    16'h535C: data_out = 8'hAF;
                    16'h535D: data_out = 8'hB0;
                    16'h535E: data_out = 8'hB1;
                    16'h535F: data_out = 8'hB2;
                    16'h5360: data_out = 8'hB3;
                    16'h5361: data_out = 8'hB4;
                    16'h5362: data_out = 8'hB5;
                    16'h5363: data_out = 8'hB6;
                    16'h5364: data_out = 8'hB7;
                    16'h5365: data_out = 8'hB8;
                    16'h5366: data_out = 8'hB9;
                    16'h5367: data_out = 8'hBA;
                    16'h5368: data_out = 8'hBB;
                    16'h5369: data_out = 8'hBC;
                    16'h536A: data_out = 8'hBD;
                    16'h536B: data_out = 8'hBE;
                    16'h536C: data_out = 8'hBF;
                    16'h536D: data_out = 8'hC0;
                    16'h536E: data_out = 8'hC1;
                    16'h536F: data_out = 8'hC2;
                    16'h5370: data_out = 8'hC3;
                    16'h5371: data_out = 8'hC4;
                    16'h5372: data_out = 8'hC5;
                    16'h5373: data_out = 8'hC6;
                    16'h5374: data_out = 8'hC7;
                    16'h5375: data_out = 8'hC8;
                    16'h5376: data_out = 8'hC9;
                    16'h5377: data_out = 8'hCA;
                    16'h5378: data_out = 8'hCB;
                    16'h5379: data_out = 8'hCC;
                    16'h537A: data_out = 8'hCD;
                    16'h537B: data_out = 8'hCE;
                    16'h537C: data_out = 8'hCF;
                    16'h537D: data_out = 8'hD0;
                    16'h537E: data_out = 8'hD1;
                    16'h537F: data_out = 8'hD2;
                    16'h5380: data_out = 8'h53;
                    16'h5381: data_out = 8'h52;
                    16'h5382: data_out = 8'h51;
                    16'h5383: data_out = 8'h50;
                    16'h5384: data_out = 8'h4F;
                    16'h5385: data_out = 8'h4E;
                    16'h5386: data_out = 8'h4D;
                    16'h5387: data_out = 8'h4C;
                    16'h5388: data_out = 8'h4B;
                    16'h5389: data_out = 8'h4A;
                    16'h538A: data_out = 8'h49;
                    16'h538B: data_out = 8'h48;
                    16'h538C: data_out = 8'h47;
                    16'h538D: data_out = 8'h46;
                    16'h538E: data_out = 8'h45;
                    16'h538F: data_out = 8'h44;
                    16'h5390: data_out = 8'h43;
                    16'h5391: data_out = 8'h42;
                    16'h5392: data_out = 8'h41;
                    16'h5393: data_out = 8'h40;
                    16'h5394: data_out = 8'h3F;
                    16'h5395: data_out = 8'h3E;
                    16'h5396: data_out = 8'h3D;
                    16'h5397: data_out = 8'h3C;
                    16'h5398: data_out = 8'h3B;
                    16'h5399: data_out = 8'h3A;
                    16'h539A: data_out = 8'h39;
                    16'h539B: data_out = 8'h38;
                    16'h539C: data_out = 8'h37;
                    16'h539D: data_out = 8'h36;
                    16'h539E: data_out = 8'h35;
                    16'h539F: data_out = 8'h34;
                    16'h53A0: data_out = 8'h33;
                    16'h53A1: data_out = 8'h32;
                    16'h53A2: data_out = 8'h31;
                    16'h53A3: data_out = 8'h30;
                    16'h53A4: data_out = 8'h2F;
                    16'h53A5: data_out = 8'h2E;
                    16'h53A6: data_out = 8'h2D;
                    16'h53A7: data_out = 8'h2C;
                    16'h53A8: data_out = 8'h2B;
                    16'h53A9: data_out = 8'h2A;
                    16'h53AA: data_out = 8'h29;
                    16'h53AB: data_out = 8'h28;
                    16'h53AC: data_out = 8'h27;
                    16'h53AD: data_out = 8'h26;
                    16'h53AE: data_out = 8'h25;
                    16'h53AF: data_out = 8'h24;
                    16'h53B0: data_out = 8'h23;
                    16'h53B1: data_out = 8'h22;
                    16'h53B2: data_out = 8'h21;
                    16'h53B3: data_out = 8'h20;
                    16'h53B4: data_out = 8'h1F;
                    16'h53B5: data_out = 8'h1E;
                    16'h53B6: data_out = 8'h1D;
                    16'h53B7: data_out = 8'h1C;
                    16'h53B8: data_out = 8'h1B;
                    16'h53B9: data_out = 8'h1A;
                    16'h53BA: data_out = 8'h19;
                    16'h53BB: data_out = 8'h18;
                    16'h53BC: data_out = 8'h17;
                    16'h53BD: data_out = 8'h16;
                    16'h53BE: data_out = 8'h15;
                    16'h53BF: data_out = 8'h14;
                    16'h53C0: data_out = 8'h13;
                    16'h53C1: data_out = 8'h12;
                    16'h53C2: data_out = 8'h11;
                    16'h53C3: data_out = 8'h10;
                    16'h53C4: data_out = 8'hF;
                    16'h53C5: data_out = 8'hE;
                    16'h53C6: data_out = 8'hD;
                    16'h53C7: data_out = 8'hC;
                    16'h53C8: data_out = 8'hB;
                    16'h53C9: data_out = 8'hA;
                    16'h53CA: data_out = 8'h9;
                    16'h53CB: data_out = 8'h8;
                    16'h53CC: data_out = 8'h7;
                    16'h53CD: data_out = 8'h6;
                    16'h53CE: data_out = 8'h5;
                    16'h53CF: data_out = 8'h4;
                    16'h53D0: data_out = 8'h3;
                    16'h53D1: data_out = 8'h2;
                    16'h53D2: data_out = 8'h1;
                    16'h53D3: data_out = 8'h0;
                    16'h53D4: data_out = 8'h81;
                    16'h53D5: data_out = 8'h82;
                    16'h53D6: data_out = 8'h83;
                    16'h53D7: data_out = 8'h84;
                    16'h53D8: data_out = 8'h85;
                    16'h53D9: data_out = 8'h86;
                    16'h53DA: data_out = 8'h87;
                    16'h53DB: data_out = 8'h88;
                    16'h53DC: data_out = 8'h89;
                    16'h53DD: data_out = 8'h8A;
                    16'h53DE: data_out = 8'h8B;
                    16'h53DF: data_out = 8'h8C;
                    16'h53E0: data_out = 8'h8D;
                    16'h53E1: data_out = 8'h8E;
                    16'h53E2: data_out = 8'h8F;
                    16'h53E3: data_out = 8'h90;
                    16'h53E4: data_out = 8'h91;
                    16'h53E5: data_out = 8'h92;
                    16'h53E6: data_out = 8'h93;
                    16'h53E7: data_out = 8'h94;
                    16'h53E8: data_out = 8'h95;
                    16'h53E9: data_out = 8'h96;
                    16'h53EA: data_out = 8'h97;
                    16'h53EB: data_out = 8'h98;
                    16'h53EC: data_out = 8'h99;
                    16'h53ED: data_out = 8'h9A;
                    16'h53EE: data_out = 8'h9B;
                    16'h53EF: data_out = 8'h9C;
                    16'h53F0: data_out = 8'h9D;
                    16'h53F1: data_out = 8'h9E;
                    16'h53F2: data_out = 8'h9F;
                    16'h53F3: data_out = 8'hA0;
                    16'h53F4: data_out = 8'hA1;
                    16'h53F5: data_out = 8'hA2;
                    16'h53F6: data_out = 8'hA3;
                    16'h53F7: data_out = 8'hA4;
                    16'h53F8: data_out = 8'hA5;
                    16'h53F9: data_out = 8'hA6;
                    16'h53FA: data_out = 8'hA7;
                    16'h53FB: data_out = 8'hA8;
                    16'h53FC: data_out = 8'hA9;
                    16'h53FD: data_out = 8'hAA;
                    16'h53FE: data_out = 8'hAB;
                    16'h53FF: data_out = 8'hAC;
                    16'h5400: data_out = 8'h54;
                    16'h5401: data_out = 8'h55;
                    16'h5402: data_out = 8'h56;
                    16'h5403: data_out = 8'h57;
                    16'h5404: data_out = 8'h58;
                    16'h5405: data_out = 8'h59;
                    16'h5406: data_out = 8'h5A;
                    16'h5407: data_out = 8'h5B;
                    16'h5408: data_out = 8'h5C;
                    16'h5409: data_out = 8'h5D;
                    16'h540A: data_out = 8'h5E;
                    16'h540B: data_out = 8'h5F;
                    16'h540C: data_out = 8'h60;
                    16'h540D: data_out = 8'h61;
                    16'h540E: data_out = 8'h62;
                    16'h540F: data_out = 8'h63;
                    16'h5410: data_out = 8'h64;
                    16'h5411: data_out = 8'h65;
                    16'h5412: data_out = 8'h66;
                    16'h5413: data_out = 8'h67;
                    16'h5414: data_out = 8'h68;
                    16'h5415: data_out = 8'h69;
                    16'h5416: data_out = 8'h6A;
                    16'h5417: data_out = 8'h6B;
                    16'h5418: data_out = 8'h6C;
                    16'h5419: data_out = 8'h6D;
                    16'h541A: data_out = 8'h6E;
                    16'h541B: data_out = 8'h6F;
                    16'h541C: data_out = 8'h70;
                    16'h541D: data_out = 8'h71;
                    16'h541E: data_out = 8'h72;
                    16'h541F: data_out = 8'h73;
                    16'h5420: data_out = 8'h74;
                    16'h5421: data_out = 8'h75;
                    16'h5422: data_out = 8'h76;
                    16'h5423: data_out = 8'h77;
                    16'h5424: data_out = 8'h78;
                    16'h5425: data_out = 8'h79;
                    16'h5426: data_out = 8'h7A;
                    16'h5427: data_out = 8'h7B;
                    16'h5428: data_out = 8'h7C;
                    16'h5429: data_out = 8'h7D;
                    16'h542A: data_out = 8'h7E;
                    16'h542B: data_out = 8'h7F;
                    16'h542C: data_out = 8'h80;
                    16'h542D: data_out = 8'h81;
                    16'h542E: data_out = 8'h82;
                    16'h542F: data_out = 8'h83;
                    16'h5430: data_out = 8'h84;
                    16'h5431: data_out = 8'h85;
                    16'h5432: data_out = 8'h86;
                    16'h5433: data_out = 8'h87;
                    16'h5434: data_out = 8'h88;
                    16'h5435: data_out = 8'h89;
                    16'h5436: data_out = 8'h8A;
                    16'h5437: data_out = 8'h8B;
                    16'h5438: data_out = 8'h8C;
                    16'h5439: data_out = 8'h8D;
                    16'h543A: data_out = 8'h8E;
                    16'h543B: data_out = 8'h8F;
                    16'h543C: data_out = 8'h90;
                    16'h543D: data_out = 8'h91;
                    16'h543E: data_out = 8'h92;
                    16'h543F: data_out = 8'h93;
                    16'h5440: data_out = 8'h94;
                    16'h5441: data_out = 8'h95;
                    16'h5442: data_out = 8'h96;
                    16'h5443: data_out = 8'h97;
                    16'h5444: data_out = 8'h98;
                    16'h5445: data_out = 8'h99;
                    16'h5446: data_out = 8'h9A;
                    16'h5447: data_out = 8'h9B;
                    16'h5448: data_out = 8'h9C;
                    16'h5449: data_out = 8'h9D;
                    16'h544A: data_out = 8'h9E;
                    16'h544B: data_out = 8'h9F;
                    16'h544C: data_out = 8'hA0;
                    16'h544D: data_out = 8'hA1;
                    16'h544E: data_out = 8'hA2;
                    16'h544F: data_out = 8'hA3;
                    16'h5450: data_out = 8'hA4;
                    16'h5451: data_out = 8'hA5;
                    16'h5452: data_out = 8'hA6;
                    16'h5453: data_out = 8'hA7;
                    16'h5454: data_out = 8'hA8;
                    16'h5455: data_out = 8'hA9;
                    16'h5456: data_out = 8'hAA;
                    16'h5457: data_out = 8'hAB;
                    16'h5458: data_out = 8'hAC;
                    16'h5459: data_out = 8'hAD;
                    16'h545A: data_out = 8'hAE;
                    16'h545B: data_out = 8'hAF;
                    16'h545C: data_out = 8'hB0;
                    16'h545D: data_out = 8'hB1;
                    16'h545E: data_out = 8'hB2;
                    16'h545F: data_out = 8'hB3;
                    16'h5460: data_out = 8'hB4;
                    16'h5461: data_out = 8'hB5;
                    16'h5462: data_out = 8'hB6;
                    16'h5463: data_out = 8'hB7;
                    16'h5464: data_out = 8'hB8;
                    16'h5465: data_out = 8'hB9;
                    16'h5466: data_out = 8'hBA;
                    16'h5467: data_out = 8'hBB;
                    16'h5468: data_out = 8'hBC;
                    16'h5469: data_out = 8'hBD;
                    16'h546A: data_out = 8'hBE;
                    16'h546B: data_out = 8'hBF;
                    16'h546C: data_out = 8'hC0;
                    16'h546D: data_out = 8'hC1;
                    16'h546E: data_out = 8'hC2;
                    16'h546F: data_out = 8'hC3;
                    16'h5470: data_out = 8'hC4;
                    16'h5471: data_out = 8'hC5;
                    16'h5472: data_out = 8'hC6;
                    16'h5473: data_out = 8'hC7;
                    16'h5474: data_out = 8'hC8;
                    16'h5475: data_out = 8'hC9;
                    16'h5476: data_out = 8'hCA;
                    16'h5477: data_out = 8'hCB;
                    16'h5478: data_out = 8'hCC;
                    16'h5479: data_out = 8'hCD;
                    16'h547A: data_out = 8'hCE;
                    16'h547B: data_out = 8'hCF;
                    16'h547C: data_out = 8'hD0;
                    16'h547D: data_out = 8'hD1;
                    16'h547E: data_out = 8'hD2;
                    16'h547F: data_out = 8'hD3;
                    16'h5480: data_out = 8'h54;
                    16'h5481: data_out = 8'h53;
                    16'h5482: data_out = 8'h52;
                    16'h5483: data_out = 8'h51;
                    16'h5484: data_out = 8'h50;
                    16'h5485: data_out = 8'h4F;
                    16'h5486: data_out = 8'h4E;
                    16'h5487: data_out = 8'h4D;
                    16'h5488: data_out = 8'h4C;
                    16'h5489: data_out = 8'h4B;
                    16'h548A: data_out = 8'h4A;
                    16'h548B: data_out = 8'h49;
                    16'h548C: data_out = 8'h48;
                    16'h548D: data_out = 8'h47;
                    16'h548E: data_out = 8'h46;
                    16'h548F: data_out = 8'h45;
                    16'h5490: data_out = 8'h44;
                    16'h5491: data_out = 8'h43;
                    16'h5492: data_out = 8'h42;
                    16'h5493: data_out = 8'h41;
                    16'h5494: data_out = 8'h40;
                    16'h5495: data_out = 8'h3F;
                    16'h5496: data_out = 8'h3E;
                    16'h5497: data_out = 8'h3D;
                    16'h5498: data_out = 8'h3C;
                    16'h5499: data_out = 8'h3B;
                    16'h549A: data_out = 8'h3A;
                    16'h549B: data_out = 8'h39;
                    16'h549C: data_out = 8'h38;
                    16'h549D: data_out = 8'h37;
                    16'h549E: data_out = 8'h36;
                    16'h549F: data_out = 8'h35;
                    16'h54A0: data_out = 8'h34;
                    16'h54A1: data_out = 8'h33;
                    16'h54A2: data_out = 8'h32;
                    16'h54A3: data_out = 8'h31;
                    16'h54A4: data_out = 8'h30;
                    16'h54A5: data_out = 8'h2F;
                    16'h54A6: data_out = 8'h2E;
                    16'h54A7: data_out = 8'h2D;
                    16'h54A8: data_out = 8'h2C;
                    16'h54A9: data_out = 8'h2B;
                    16'h54AA: data_out = 8'h2A;
                    16'h54AB: data_out = 8'h29;
                    16'h54AC: data_out = 8'h28;
                    16'h54AD: data_out = 8'h27;
                    16'h54AE: data_out = 8'h26;
                    16'h54AF: data_out = 8'h25;
                    16'h54B0: data_out = 8'h24;
                    16'h54B1: data_out = 8'h23;
                    16'h54B2: data_out = 8'h22;
                    16'h54B3: data_out = 8'h21;
                    16'h54B4: data_out = 8'h20;
                    16'h54B5: data_out = 8'h1F;
                    16'h54B6: data_out = 8'h1E;
                    16'h54B7: data_out = 8'h1D;
                    16'h54B8: data_out = 8'h1C;
                    16'h54B9: data_out = 8'h1B;
                    16'h54BA: data_out = 8'h1A;
                    16'h54BB: data_out = 8'h19;
                    16'h54BC: data_out = 8'h18;
                    16'h54BD: data_out = 8'h17;
                    16'h54BE: data_out = 8'h16;
                    16'h54BF: data_out = 8'h15;
                    16'h54C0: data_out = 8'h14;
                    16'h54C1: data_out = 8'h13;
                    16'h54C2: data_out = 8'h12;
                    16'h54C3: data_out = 8'h11;
                    16'h54C4: data_out = 8'h10;
                    16'h54C5: data_out = 8'hF;
                    16'h54C6: data_out = 8'hE;
                    16'h54C7: data_out = 8'hD;
                    16'h54C8: data_out = 8'hC;
                    16'h54C9: data_out = 8'hB;
                    16'h54CA: data_out = 8'hA;
                    16'h54CB: data_out = 8'h9;
                    16'h54CC: data_out = 8'h8;
                    16'h54CD: data_out = 8'h7;
                    16'h54CE: data_out = 8'h6;
                    16'h54CF: data_out = 8'h5;
                    16'h54D0: data_out = 8'h4;
                    16'h54D1: data_out = 8'h3;
                    16'h54D2: data_out = 8'h2;
                    16'h54D3: data_out = 8'h1;
                    16'h54D4: data_out = 8'h0;
                    16'h54D5: data_out = 8'h81;
                    16'h54D6: data_out = 8'h82;
                    16'h54D7: data_out = 8'h83;
                    16'h54D8: data_out = 8'h84;
                    16'h54D9: data_out = 8'h85;
                    16'h54DA: data_out = 8'h86;
                    16'h54DB: data_out = 8'h87;
                    16'h54DC: data_out = 8'h88;
                    16'h54DD: data_out = 8'h89;
                    16'h54DE: data_out = 8'h8A;
                    16'h54DF: data_out = 8'h8B;
                    16'h54E0: data_out = 8'h8C;
                    16'h54E1: data_out = 8'h8D;
                    16'h54E2: data_out = 8'h8E;
                    16'h54E3: data_out = 8'h8F;
                    16'h54E4: data_out = 8'h90;
                    16'h54E5: data_out = 8'h91;
                    16'h54E6: data_out = 8'h92;
                    16'h54E7: data_out = 8'h93;
                    16'h54E8: data_out = 8'h94;
                    16'h54E9: data_out = 8'h95;
                    16'h54EA: data_out = 8'h96;
                    16'h54EB: data_out = 8'h97;
                    16'h54EC: data_out = 8'h98;
                    16'h54ED: data_out = 8'h99;
                    16'h54EE: data_out = 8'h9A;
                    16'h54EF: data_out = 8'h9B;
                    16'h54F0: data_out = 8'h9C;
                    16'h54F1: data_out = 8'h9D;
                    16'h54F2: data_out = 8'h9E;
                    16'h54F3: data_out = 8'h9F;
                    16'h54F4: data_out = 8'hA0;
                    16'h54F5: data_out = 8'hA1;
                    16'h54F6: data_out = 8'hA2;
                    16'h54F7: data_out = 8'hA3;
                    16'h54F8: data_out = 8'hA4;
                    16'h54F9: data_out = 8'hA5;
                    16'h54FA: data_out = 8'hA6;
                    16'h54FB: data_out = 8'hA7;
                    16'h54FC: data_out = 8'hA8;
                    16'h54FD: data_out = 8'hA9;
                    16'h54FE: data_out = 8'hAA;
                    16'h54FF: data_out = 8'hAB;
                    16'h5500: data_out = 8'h55;
                    16'h5501: data_out = 8'h56;
                    16'h5502: data_out = 8'h57;
                    16'h5503: data_out = 8'h58;
                    16'h5504: data_out = 8'h59;
                    16'h5505: data_out = 8'h5A;
                    16'h5506: data_out = 8'h5B;
                    16'h5507: data_out = 8'h5C;
                    16'h5508: data_out = 8'h5D;
                    16'h5509: data_out = 8'h5E;
                    16'h550A: data_out = 8'h5F;
                    16'h550B: data_out = 8'h60;
                    16'h550C: data_out = 8'h61;
                    16'h550D: data_out = 8'h62;
                    16'h550E: data_out = 8'h63;
                    16'h550F: data_out = 8'h64;
                    16'h5510: data_out = 8'h65;
                    16'h5511: data_out = 8'h66;
                    16'h5512: data_out = 8'h67;
                    16'h5513: data_out = 8'h68;
                    16'h5514: data_out = 8'h69;
                    16'h5515: data_out = 8'h6A;
                    16'h5516: data_out = 8'h6B;
                    16'h5517: data_out = 8'h6C;
                    16'h5518: data_out = 8'h6D;
                    16'h5519: data_out = 8'h6E;
                    16'h551A: data_out = 8'h6F;
                    16'h551B: data_out = 8'h70;
                    16'h551C: data_out = 8'h71;
                    16'h551D: data_out = 8'h72;
                    16'h551E: data_out = 8'h73;
                    16'h551F: data_out = 8'h74;
                    16'h5520: data_out = 8'h75;
                    16'h5521: data_out = 8'h76;
                    16'h5522: data_out = 8'h77;
                    16'h5523: data_out = 8'h78;
                    16'h5524: data_out = 8'h79;
                    16'h5525: data_out = 8'h7A;
                    16'h5526: data_out = 8'h7B;
                    16'h5527: data_out = 8'h7C;
                    16'h5528: data_out = 8'h7D;
                    16'h5529: data_out = 8'h7E;
                    16'h552A: data_out = 8'h7F;
                    16'h552B: data_out = 8'h80;
                    16'h552C: data_out = 8'h81;
                    16'h552D: data_out = 8'h82;
                    16'h552E: data_out = 8'h83;
                    16'h552F: data_out = 8'h84;
                    16'h5530: data_out = 8'h85;
                    16'h5531: data_out = 8'h86;
                    16'h5532: data_out = 8'h87;
                    16'h5533: data_out = 8'h88;
                    16'h5534: data_out = 8'h89;
                    16'h5535: data_out = 8'h8A;
                    16'h5536: data_out = 8'h8B;
                    16'h5537: data_out = 8'h8C;
                    16'h5538: data_out = 8'h8D;
                    16'h5539: data_out = 8'h8E;
                    16'h553A: data_out = 8'h8F;
                    16'h553B: data_out = 8'h90;
                    16'h553C: data_out = 8'h91;
                    16'h553D: data_out = 8'h92;
                    16'h553E: data_out = 8'h93;
                    16'h553F: data_out = 8'h94;
                    16'h5540: data_out = 8'h95;
                    16'h5541: data_out = 8'h96;
                    16'h5542: data_out = 8'h97;
                    16'h5543: data_out = 8'h98;
                    16'h5544: data_out = 8'h99;
                    16'h5545: data_out = 8'h9A;
                    16'h5546: data_out = 8'h9B;
                    16'h5547: data_out = 8'h9C;
                    16'h5548: data_out = 8'h9D;
                    16'h5549: data_out = 8'h9E;
                    16'h554A: data_out = 8'h9F;
                    16'h554B: data_out = 8'hA0;
                    16'h554C: data_out = 8'hA1;
                    16'h554D: data_out = 8'hA2;
                    16'h554E: data_out = 8'hA3;
                    16'h554F: data_out = 8'hA4;
                    16'h5550: data_out = 8'hA5;
                    16'h5551: data_out = 8'hA6;
                    16'h5552: data_out = 8'hA7;
                    16'h5553: data_out = 8'hA8;
                    16'h5554: data_out = 8'hA9;
                    16'h5555: data_out = 8'hAA;
                    16'h5556: data_out = 8'hAB;
                    16'h5557: data_out = 8'hAC;
                    16'h5558: data_out = 8'hAD;
                    16'h5559: data_out = 8'hAE;
                    16'h555A: data_out = 8'hAF;
                    16'h555B: data_out = 8'hB0;
                    16'h555C: data_out = 8'hB1;
                    16'h555D: data_out = 8'hB2;
                    16'h555E: data_out = 8'hB3;
                    16'h555F: data_out = 8'hB4;
                    16'h5560: data_out = 8'hB5;
                    16'h5561: data_out = 8'hB6;
                    16'h5562: data_out = 8'hB7;
                    16'h5563: data_out = 8'hB8;
                    16'h5564: data_out = 8'hB9;
                    16'h5565: data_out = 8'hBA;
                    16'h5566: data_out = 8'hBB;
                    16'h5567: data_out = 8'hBC;
                    16'h5568: data_out = 8'hBD;
                    16'h5569: data_out = 8'hBE;
                    16'h556A: data_out = 8'hBF;
                    16'h556B: data_out = 8'hC0;
                    16'h556C: data_out = 8'hC1;
                    16'h556D: data_out = 8'hC2;
                    16'h556E: data_out = 8'hC3;
                    16'h556F: data_out = 8'hC4;
                    16'h5570: data_out = 8'hC5;
                    16'h5571: data_out = 8'hC6;
                    16'h5572: data_out = 8'hC7;
                    16'h5573: data_out = 8'hC8;
                    16'h5574: data_out = 8'hC9;
                    16'h5575: data_out = 8'hCA;
                    16'h5576: data_out = 8'hCB;
                    16'h5577: data_out = 8'hCC;
                    16'h5578: data_out = 8'hCD;
                    16'h5579: data_out = 8'hCE;
                    16'h557A: data_out = 8'hCF;
                    16'h557B: data_out = 8'hD0;
                    16'h557C: data_out = 8'hD1;
                    16'h557D: data_out = 8'hD2;
                    16'h557E: data_out = 8'hD3;
                    16'h557F: data_out = 8'hD4;
                    16'h5580: data_out = 8'h55;
                    16'h5581: data_out = 8'h54;
                    16'h5582: data_out = 8'h53;
                    16'h5583: data_out = 8'h52;
                    16'h5584: data_out = 8'h51;
                    16'h5585: data_out = 8'h50;
                    16'h5586: data_out = 8'h4F;
                    16'h5587: data_out = 8'h4E;
                    16'h5588: data_out = 8'h4D;
                    16'h5589: data_out = 8'h4C;
                    16'h558A: data_out = 8'h4B;
                    16'h558B: data_out = 8'h4A;
                    16'h558C: data_out = 8'h49;
                    16'h558D: data_out = 8'h48;
                    16'h558E: data_out = 8'h47;
                    16'h558F: data_out = 8'h46;
                    16'h5590: data_out = 8'h45;
                    16'h5591: data_out = 8'h44;
                    16'h5592: data_out = 8'h43;
                    16'h5593: data_out = 8'h42;
                    16'h5594: data_out = 8'h41;
                    16'h5595: data_out = 8'h40;
                    16'h5596: data_out = 8'h3F;
                    16'h5597: data_out = 8'h3E;
                    16'h5598: data_out = 8'h3D;
                    16'h5599: data_out = 8'h3C;
                    16'h559A: data_out = 8'h3B;
                    16'h559B: data_out = 8'h3A;
                    16'h559C: data_out = 8'h39;
                    16'h559D: data_out = 8'h38;
                    16'h559E: data_out = 8'h37;
                    16'h559F: data_out = 8'h36;
                    16'h55A0: data_out = 8'h35;
                    16'h55A1: data_out = 8'h34;
                    16'h55A2: data_out = 8'h33;
                    16'h55A3: data_out = 8'h32;
                    16'h55A4: data_out = 8'h31;
                    16'h55A5: data_out = 8'h30;
                    16'h55A6: data_out = 8'h2F;
                    16'h55A7: data_out = 8'h2E;
                    16'h55A8: data_out = 8'h2D;
                    16'h55A9: data_out = 8'h2C;
                    16'h55AA: data_out = 8'h2B;
                    16'h55AB: data_out = 8'h2A;
                    16'h55AC: data_out = 8'h29;
                    16'h55AD: data_out = 8'h28;
                    16'h55AE: data_out = 8'h27;
                    16'h55AF: data_out = 8'h26;
                    16'h55B0: data_out = 8'h25;
                    16'h55B1: data_out = 8'h24;
                    16'h55B2: data_out = 8'h23;
                    16'h55B3: data_out = 8'h22;
                    16'h55B4: data_out = 8'h21;
                    16'h55B5: data_out = 8'h20;
                    16'h55B6: data_out = 8'h1F;
                    16'h55B7: data_out = 8'h1E;
                    16'h55B8: data_out = 8'h1D;
                    16'h55B9: data_out = 8'h1C;
                    16'h55BA: data_out = 8'h1B;
                    16'h55BB: data_out = 8'h1A;
                    16'h55BC: data_out = 8'h19;
                    16'h55BD: data_out = 8'h18;
                    16'h55BE: data_out = 8'h17;
                    16'h55BF: data_out = 8'h16;
                    16'h55C0: data_out = 8'h15;
                    16'h55C1: data_out = 8'h14;
                    16'h55C2: data_out = 8'h13;
                    16'h55C3: data_out = 8'h12;
                    16'h55C4: data_out = 8'h11;
                    16'h55C5: data_out = 8'h10;
                    16'h55C6: data_out = 8'hF;
                    16'h55C7: data_out = 8'hE;
                    16'h55C8: data_out = 8'hD;
                    16'h55C9: data_out = 8'hC;
                    16'h55CA: data_out = 8'hB;
                    16'h55CB: data_out = 8'hA;
                    16'h55CC: data_out = 8'h9;
                    16'h55CD: data_out = 8'h8;
                    16'h55CE: data_out = 8'h7;
                    16'h55CF: data_out = 8'h6;
                    16'h55D0: data_out = 8'h5;
                    16'h55D1: data_out = 8'h4;
                    16'h55D2: data_out = 8'h3;
                    16'h55D3: data_out = 8'h2;
                    16'h55D4: data_out = 8'h1;
                    16'h55D5: data_out = 8'h0;
                    16'h55D6: data_out = 8'h81;
                    16'h55D7: data_out = 8'h82;
                    16'h55D8: data_out = 8'h83;
                    16'h55D9: data_out = 8'h84;
                    16'h55DA: data_out = 8'h85;
                    16'h55DB: data_out = 8'h86;
                    16'h55DC: data_out = 8'h87;
                    16'h55DD: data_out = 8'h88;
                    16'h55DE: data_out = 8'h89;
                    16'h55DF: data_out = 8'h8A;
                    16'h55E0: data_out = 8'h8B;
                    16'h55E1: data_out = 8'h8C;
                    16'h55E2: data_out = 8'h8D;
                    16'h55E3: data_out = 8'h8E;
                    16'h55E4: data_out = 8'h8F;
                    16'h55E5: data_out = 8'h90;
                    16'h55E6: data_out = 8'h91;
                    16'h55E7: data_out = 8'h92;
                    16'h55E8: data_out = 8'h93;
                    16'h55E9: data_out = 8'h94;
                    16'h55EA: data_out = 8'h95;
                    16'h55EB: data_out = 8'h96;
                    16'h55EC: data_out = 8'h97;
                    16'h55ED: data_out = 8'h98;
                    16'h55EE: data_out = 8'h99;
                    16'h55EF: data_out = 8'h9A;
                    16'h55F0: data_out = 8'h9B;
                    16'h55F1: data_out = 8'h9C;
                    16'h55F2: data_out = 8'h9D;
                    16'h55F3: data_out = 8'h9E;
                    16'h55F4: data_out = 8'h9F;
                    16'h55F5: data_out = 8'hA0;
                    16'h55F6: data_out = 8'hA1;
                    16'h55F7: data_out = 8'hA2;
                    16'h55F8: data_out = 8'hA3;
                    16'h55F9: data_out = 8'hA4;
                    16'h55FA: data_out = 8'hA5;
                    16'h55FB: data_out = 8'hA6;
                    16'h55FC: data_out = 8'hA7;
                    16'h55FD: data_out = 8'hA8;
                    16'h55FE: data_out = 8'hA9;
                    16'h55FF: data_out = 8'hAA;
                    16'h5600: data_out = 8'h56;
                    16'h5601: data_out = 8'h57;
                    16'h5602: data_out = 8'h58;
                    16'h5603: data_out = 8'h59;
                    16'h5604: data_out = 8'h5A;
                    16'h5605: data_out = 8'h5B;
                    16'h5606: data_out = 8'h5C;
                    16'h5607: data_out = 8'h5D;
                    16'h5608: data_out = 8'h5E;
                    16'h5609: data_out = 8'h5F;
                    16'h560A: data_out = 8'h60;
                    16'h560B: data_out = 8'h61;
                    16'h560C: data_out = 8'h62;
                    16'h560D: data_out = 8'h63;
                    16'h560E: data_out = 8'h64;
                    16'h560F: data_out = 8'h65;
                    16'h5610: data_out = 8'h66;
                    16'h5611: data_out = 8'h67;
                    16'h5612: data_out = 8'h68;
                    16'h5613: data_out = 8'h69;
                    16'h5614: data_out = 8'h6A;
                    16'h5615: data_out = 8'h6B;
                    16'h5616: data_out = 8'h6C;
                    16'h5617: data_out = 8'h6D;
                    16'h5618: data_out = 8'h6E;
                    16'h5619: data_out = 8'h6F;
                    16'h561A: data_out = 8'h70;
                    16'h561B: data_out = 8'h71;
                    16'h561C: data_out = 8'h72;
                    16'h561D: data_out = 8'h73;
                    16'h561E: data_out = 8'h74;
                    16'h561F: data_out = 8'h75;
                    16'h5620: data_out = 8'h76;
                    16'h5621: data_out = 8'h77;
                    16'h5622: data_out = 8'h78;
                    16'h5623: data_out = 8'h79;
                    16'h5624: data_out = 8'h7A;
                    16'h5625: data_out = 8'h7B;
                    16'h5626: data_out = 8'h7C;
                    16'h5627: data_out = 8'h7D;
                    16'h5628: data_out = 8'h7E;
                    16'h5629: data_out = 8'h7F;
                    16'h562A: data_out = 8'h80;
                    16'h562B: data_out = 8'h81;
                    16'h562C: data_out = 8'h82;
                    16'h562D: data_out = 8'h83;
                    16'h562E: data_out = 8'h84;
                    16'h562F: data_out = 8'h85;
                    16'h5630: data_out = 8'h86;
                    16'h5631: data_out = 8'h87;
                    16'h5632: data_out = 8'h88;
                    16'h5633: data_out = 8'h89;
                    16'h5634: data_out = 8'h8A;
                    16'h5635: data_out = 8'h8B;
                    16'h5636: data_out = 8'h8C;
                    16'h5637: data_out = 8'h8D;
                    16'h5638: data_out = 8'h8E;
                    16'h5639: data_out = 8'h8F;
                    16'h563A: data_out = 8'h90;
                    16'h563B: data_out = 8'h91;
                    16'h563C: data_out = 8'h92;
                    16'h563D: data_out = 8'h93;
                    16'h563E: data_out = 8'h94;
                    16'h563F: data_out = 8'h95;
                    16'h5640: data_out = 8'h96;
                    16'h5641: data_out = 8'h97;
                    16'h5642: data_out = 8'h98;
                    16'h5643: data_out = 8'h99;
                    16'h5644: data_out = 8'h9A;
                    16'h5645: data_out = 8'h9B;
                    16'h5646: data_out = 8'h9C;
                    16'h5647: data_out = 8'h9D;
                    16'h5648: data_out = 8'h9E;
                    16'h5649: data_out = 8'h9F;
                    16'h564A: data_out = 8'hA0;
                    16'h564B: data_out = 8'hA1;
                    16'h564C: data_out = 8'hA2;
                    16'h564D: data_out = 8'hA3;
                    16'h564E: data_out = 8'hA4;
                    16'h564F: data_out = 8'hA5;
                    16'h5650: data_out = 8'hA6;
                    16'h5651: data_out = 8'hA7;
                    16'h5652: data_out = 8'hA8;
                    16'h5653: data_out = 8'hA9;
                    16'h5654: data_out = 8'hAA;
                    16'h5655: data_out = 8'hAB;
                    16'h5656: data_out = 8'hAC;
                    16'h5657: data_out = 8'hAD;
                    16'h5658: data_out = 8'hAE;
                    16'h5659: data_out = 8'hAF;
                    16'h565A: data_out = 8'hB0;
                    16'h565B: data_out = 8'hB1;
                    16'h565C: data_out = 8'hB2;
                    16'h565D: data_out = 8'hB3;
                    16'h565E: data_out = 8'hB4;
                    16'h565F: data_out = 8'hB5;
                    16'h5660: data_out = 8'hB6;
                    16'h5661: data_out = 8'hB7;
                    16'h5662: data_out = 8'hB8;
                    16'h5663: data_out = 8'hB9;
                    16'h5664: data_out = 8'hBA;
                    16'h5665: data_out = 8'hBB;
                    16'h5666: data_out = 8'hBC;
                    16'h5667: data_out = 8'hBD;
                    16'h5668: data_out = 8'hBE;
                    16'h5669: data_out = 8'hBF;
                    16'h566A: data_out = 8'hC0;
                    16'h566B: data_out = 8'hC1;
                    16'h566C: data_out = 8'hC2;
                    16'h566D: data_out = 8'hC3;
                    16'h566E: data_out = 8'hC4;
                    16'h566F: data_out = 8'hC5;
                    16'h5670: data_out = 8'hC6;
                    16'h5671: data_out = 8'hC7;
                    16'h5672: data_out = 8'hC8;
                    16'h5673: data_out = 8'hC9;
                    16'h5674: data_out = 8'hCA;
                    16'h5675: data_out = 8'hCB;
                    16'h5676: data_out = 8'hCC;
                    16'h5677: data_out = 8'hCD;
                    16'h5678: data_out = 8'hCE;
                    16'h5679: data_out = 8'hCF;
                    16'h567A: data_out = 8'hD0;
                    16'h567B: data_out = 8'hD1;
                    16'h567C: data_out = 8'hD2;
                    16'h567D: data_out = 8'hD3;
                    16'h567E: data_out = 8'hD4;
                    16'h567F: data_out = 8'hD5;
                    16'h5680: data_out = 8'h56;
                    16'h5681: data_out = 8'h55;
                    16'h5682: data_out = 8'h54;
                    16'h5683: data_out = 8'h53;
                    16'h5684: data_out = 8'h52;
                    16'h5685: data_out = 8'h51;
                    16'h5686: data_out = 8'h50;
                    16'h5687: data_out = 8'h4F;
                    16'h5688: data_out = 8'h4E;
                    16'h5689: data_out = 8'h4D;
                    16'h568A: data_out = 8'h4C;
                    16'h568B: data_out = 8'h4B;
                    16'h568C: data_out = 8'h4A;
                    16'h568D: data_out = 8'h49;
                    16'h568E: data_out = 8'h48;
                    16'h568F: data_out = 8'h47;
                    16'h5690: data_out = 8'h46;
                    16'h5691: data_out = 8'h45;
                    16'h5692: data_out = 8'h44;
                    16'h5693: data_out = 8'h43;
                    16'h5694: data_out = 8'h42;
                    16'h5695: data_out = 8'h41;
                    16'h5696: data_out = 8'h40;
                    16'h5697: data_out = 8'h3F;
                    16'h5698: data_out = 8'h3E;
                    16'h5699: data_out = 8'h3D;
                    16'h569A: data_out = 8'h3C;
                    16'h569B: data_out = 8'h3B;
                    16'h569C: data_out = 8'h3A;
                    16'h569D: data_out = 8'h39;
                    16'h569E: data_out = 8'h38;
                    16'h569F: data_out = 8'h37;
                    16'h56A0: data_out = 8'h36;
                    16'h56A1: data_out = 8'h35;
                    16'h56A2: data_out = 8'h34;
                    16'h56A3: data_out = 8'h33;
                    16'h56A4: data_out = 8'h32;
                    16'h56A5: data_out = 8'h31;
                    16'h56A6: data_out = 8'h30;
                    16'h56A7: data_out = 8'h2F;
                    16'h56A8: data_out = 8'h2E;
                    16'h56A9: data_out = 8'h2D;
                    16'h56AA: data_out = 8'h2C;
                    16'h56AB: data_out = 8'h2B;
                    16'h56AC: data_out = 8'h2A;
                    16'h56AD: data_out = 8'h29;
                    16'h56AE: data_out = 8'h28;
                    16'h56AF: data_out = 8'h27;
                    16'h56B0: data_out = 8'h26;
                    16'h56B1: data_out = 8'h25;
                    16'h56B2: data_out = 8'h24;
                    16'h56B3: data_out = 8'h23;
                    16'h56B4: data_out = 8'h22;
                    16'h56B5: data_out = 8'h21;
                    16'h56B6: data_out = 8'h20;
                    16'h56B7: data_out = 8'h1F;
                    16'h56B8: data_out = 8'h1E;
                    16'h56B9: data_out = 8'h1D;
                    16'h56BA: data_out = 8'h1C;
                    16'h56BB: data_out = 8'h1B;
                    16'h56BC: data_out = 8'h1A;
                    16'h56BD: data_out = 8'h19;
                    16'h56BE: data_out = 8'h18;
                    16'h56BF: data_out = 8'h17;
                    16'h56C0: data_out = 8'h16;
                    16'h56C1: data_out = 8'h15;
                    16'h56C2: data_out = 8'h14;
                    16'h56C3: data_out = 8'h13;
                    16'h56C4: data_out = 8'h12;
                    16'h56C5: data_out = 8'h11;
                    16'h56C6: data_out = 8'h10;
                    16'h56C7: data_out = 8'hF;
                    16'h56C8: data_out = 8'hE;
                    16'h56C9: data_out = 8'hD;
                    16'h56CA: data_out = 8'hC;
                    16'h56CB: data_out = 8'hB;
                    16'h56CC: data_out = 8'hA;
                    16'h56CD: data_out = 8'h9;
                    16'h56CE: data_out = 8'h8;
                    16'h56CF: data_out = 8'h7;
                    16'h56D0: data_out = 8'h6;
                    16'h56D1: data_out = 8'h5;
                    16'h56D2: data_out = 8'h4;
                    16'h56D3: data_out = 8'h3;
                    16'h56D4: data_out = 8'h2;
                    16'h56D5: data_out = 8'h1;
                    16'h56D6: data_out = 8'h0;
                    16'h56D7: data_out = 8'h81;
                    16'h56D8: data_out = 8'h82;
                    16'h56D9: data_out = 8'h83;
                    16'h56DA: data_out = 8'h84;
                    16'h56DB: data_out = 8'h85;
                    16'h56DC: data_out = 8'h86;
                    16'h56DD: data_out = 8'h87;
                    16'h56DE: data_out = 8'h88;
                    16'h56DF: data_out = 8'h89;
                    16'h56E0: data_out = 8'h8A;
                    16'h56E1: data_out = 8'h8B;
                    16'h56E2: data_out = 8'h8C;
                    16'h56E3: data_out = 8'h8D;
                    16'h56E4: data_out = 8'h8E;
                    16'h56E5: data_out = 8'h8F;
                    16'h56E6: data_out = 8'h90;
                    16'h56E7: data_out = 8'h91;
                    16'h56E8: data_out = 8'h92;
                    16'h56E9: data_out = 8'h93;
                    16'h56EA: data_out = 8'h94;
                    16'h56EB: data_out = 8'h95;
                    16'h56EC: data_out = 8'h96;
                    16'h56ED: data_out = 8'h97;
                    16'h56EE: data_out = 8'h98;
                    16'h56EF: data_out = 8'h99;
                    16'h56F0: data_out = 8'h9A;
                    16'h56F1: data_out = 8'h9B;
                    16'h56F2: data_out = 8'h9C;
                    16'h56F3: data_out = 8'h9D;
                    16'h56F4: data_out = 8'h9E;
                    16'h56F5: data_out = 8'h9F;
                    16'h56F6: data_out = 8'hA0;
                    16'h56F7: data_out = 8'hA1;
                    16'h56F8: data_out = 8'hA2;
                    16'h56F9: data_out = 8'hA3;
                    16'h56FA: data_out = 8'hA4;
                    16'h56FB: data_out = 8'hA5;
                    16'h56FC: data_out = 8'hA6;
                    16'h56FD: data_out = 8'hA7;
                    16'h56FE: data_out = 8'hA8;
                    16'h56FF: data_out = 8'hA9;
                    16'h5700: data_out = 8'h57;
                    16'h5701: data_out = 8'h58;
                    16'h5702: data_out = 8'h59;
                    16'h5703: data_out = 8'h5A;
                    16'h5704: data_out = 8'h5B;
                    16'h5705: data_out = 8'h5C;
                    16'h5706: data_out = 8'h5D;
                    16'h5707: data_out = 8'h5E;
                    16'h5708: data_out = 8'h5F;
                    16'h5709: data_out = 8'h60;
                    16'h570A: data_out = 8'h61;
                    16'h570B: data_out = 8'h62;
                    16'h570C: data_out = 8'h63;
                    16'h570D: data_out = 8'h64;
                    16'h570E: data_out = 8'h65;
                    16'h570F: data_out = 8'h66;
                    16'h5710: data_out = 8'h67;
                    16'h5711: data_out = 8'h68;
                    16'h5712: data_out = 8'h69;
                    16'h5713: data_out = 8'h6A;
                    16'h5714: data_out = 8'h6B;
                    16'h5715: data_out = 8'h6C;
                    16'h5716: data_out = 8'h6D;
                    16'h5717: data_out = 8'h6E;
                    16'h5718: data_out = 8'h6F;
                    16'h5719: data_out = 8'h70;
                    16'h571A: data_out = 8'h71;
                    16'h571B: data_out = 8'h72;
                    16'h571C: data_out = 8'h73;
                    16'h571D: data_out = 8'h74;
                    16'h571E: data_out = 8'h75;
                    16'h571F: data_out = 8'h76;
                    16'h5720: data_out = 8'h77;
                    16'h5721: data_out = 8'h78;
                    16'h5722: data_out = 8'h79;
                    16'h5723: data_out = 8'h7A;
                    16'h5724: data_out = 8'h7B;
                    16'h5725: data_out = 8'h7C;
                    16'h5726: data_out = 8'h7D;
                    16'h5727: data_out = 8'h7E;
                    16'h5728: data_out = 8'h7F;
                    16'h5729: data_out = 8'h80;
                    16'h572A: data_out = 8'h81;
                    16'h572B: data_out = 8'h82;
                    16'h572C: data_out = 8'h83;
                    16'h572D: data_out = 8'h84;
                    16'h572E: data_out = 8'h85;
                    16'h572F: data_out = 8'h86;
                    16'h5730: data_out = 8'h87;
                    16'h5731: data_out = 8'h88;
                    16'h5732: data_out = 8'h89;
                    16'h5733: data_out = 8'h8A;
                    16'h5734: data_out = 8'h8B;
                    16'h5735: data_out = 8'h8C;
                    16'h5736: data_out = 8'h8D;
                    16'h5737: data_out = 8'h8E;
                    16'h5738: data_out = 8'h8F;
                    16'h5739: data_out = 8'h90;
                    16'h573A: data_out = 8'h91;
                    16'h573B: data_out = 8'h92;
                    16'h573C: data_out = 8'h93;
                    16'h573D: data_out = 8'h94;
                    16'h573E: data_out = 8'h95;
                    16'h573F: data_out = 8'h96;
                    16'h5740: data_out = 8'h97;
                    16'h5741: data_out = 8'h98;
                    16'h5742: data_out = 8'h99;
                    16'h5743: data_out = 8'h9A;
                    16'h5744: data_out = 8'h9B;
                    16'h5745: data_out = 8'h9C;
                    16'h5746: data_out = 8'h9D;
                    16'h5747: data_out = 8'h9E;
                    16'h5748: data_out = 8'h9F;
                    16'h5749: data_out = 8'hA0;
                    16'h574A: data_out = 8'hA1;
                    16'h574B: data_out = 8'hA2;
                    16'h574C: data_out = 8'hA3;
                    16'h574D: data_out = 8'hA4;
                    16'h574E: data_out = 8'hA5;
                    16'h574F: data_out = 8'hA6;
                    16'h5750: data_out = 8'hA7;
                    16'h5751: data_out = 8'hA8;
                    16'h5752: data_out = 8'hA9;
                    16'h5753: data_out = 8'hAA;
                    16'h5754: data_out = 8'hAB;
                    16'h5755: data_out = 8'hAC;
                    16'h5756: data_out = 8'hAD;
                    16'h5757: data_out = 8'hAE;
                    16'h5758: data_out = 8'hAF;
                    16'h5759: data_out = 8'hB0;
                    16'h575A: data_out = 8'hB1;
                    16'h575B: data_out = 8'hB2;
                    16'h575C: data_out = 8'hB3;
                    16'h575D: data_out = 8'hB4;
                    16'h575E: data_out = 8'hB5;
                    16'h575F: data_out = 8'hB6;
                    16'h5760: data_out = 8'hB7;
                    16'h5761: data_out = 8'hB8;
                    16'h5762: data_out = 8'hB9;
                    16'h5763: data_out = 8'hBA;
                    16'h5764: data_out = 8'hBB;
                    16'h5765: data_out = 8'hBC;
                    16'h5766: data_out = 8'hBD;
                    16'h5767: data_out = 8'hBE;
                    16'h5768: data_out = 8'hBF;
                    16'h5769: data_out = 8'hC0;
                    16'h576A: data_out = 8'hC1;
                    16'h576B: data_out = 8'hC2;
                    16'h576C: data_out = 8'hC3;
                    16'h576D: data_out = 8'hC4;
                    16'h576E: data_out = 8'hC5;
                    16'h576F: data_out = 8'hC6;
                    16'h5770: data_out = 8'hC7;
                    16'h5771: data_out = 8'hC8;
                    16'h5772: data_out = 8'hC9;
                    16'h5773: data_out = 8'hCA;
                    16'h5774: data_out = 8'hCB;
                    16'h5775: data_out = 8'hCC;
                    16'h5776: data_out = 8'hCD;
                    16'h5777: data_out = 8'hCE;
                    16'h5778: data_out = 8'hCF;
                    16'h5779: data_out = 8'hD0;
                    16'h577A: data_out = 8'hD1;
                    16'h577B: data_out = 8'hD2;
                    16'h577C: data_out = 8'hD3;
                    16'h577D: data_out = 8'hD4;
                    16'h577E: data_out = 8'hD5;
                    16'h577F: data_out = 8'hD6;
                    16'h5780: data_out = 8'h57;
                    16'h5781: data_out = 8'h56;
                    16'h5782: data_out = 8'h55;
                    16'h5783: data_out = 8'h54;
                    16'h5784: data_out = 8'h53;
                    16'h5785: data_out = 8'h52;
                    16'h5786: data_out = 8'h51;
                    16'h5787: data_out = 8'h50;
                    16'h5788: data_out = 8'h4F;
                    16'h5789: data_out = 8'h4E;
                    16'h578A: data_out = 8'h4D;
                    16'h578B: data_out = 8'h4C;
                    16'h578C: data_out = 8'h4B;
                    16'h578D: data_out = 8'h4A;
                    16'h578E: data_out = 8'h49;
                    16'h578F: data_out = 8'h48;
                    16'h5790: data_out = 8'h47;
                    16'h5791: data_out = 8'h46;
                    16'h5792: data_out = 8'h45;
                    16'h5793: data_out = 8'h44;
                    16'h5794: data_out = 8'h43;
                    16'h5795: data_out = 8'h42;
                    16'h5796: data_out = 8'h41;
                    16'h5797: data_out = 8'h40;
                    16'h5798: data_out = 8'h3F;
                    16'h5799: data_out = 8'h3E;
                    16'h579A: data_out = 8'h3D;
                    16'h579B: data_out = 8'h3C;
                    16'h579C: data_out = 8'h3B;
                    16'h579D: data_out = 8'h3A;
                    16'h579E: data_out = 8'h39;
                    16'h579F: data_out = 8'h38;
                    16'h57A0: data_out = 8'h37;
                    16'h57A1: data_out = 8'h36;
                    16'h57A2: data_out = 8'h35;
                    16'h57A3: data_out = 8'h34;
                    16'h57A4: data_out = 8'h33;
                    16'h57A5: data_out = 8'h32;
                    16'h57A6: data_out = 8'h31;
                    16'h57A7: data_out = 8'h30;
                    16'h57A8: data_out = 8'h2F;
                    16'h57A9: data_out = 8'h2E;
                    16'h57AA: data_out = 8'h2D;
                    16'h57AB: data_out = 8'h2C;
                    16'h57AC: data_out = 8'h2B;
                    16'h57AD: data_out = 8'h2A;
                    16'h57AE: data_out = 8'h29;
                    16'h57AF: data_out = 8'h28;
                    16'h57B0: data_out = 8'h27;
                    16'h57B1: data_out = 8'h26;
                    16'h57B2: data_out = 8'h25;
                    16'h57B3: data_out = 8'h24;
                    16'h57B4: data_out = 8'h23;
                    16'h57B5: data_out = 8'h22;
                    16'h57B6: data_out = 8'h21;
                    16'h57B7: data_out = 8'h20;
                    16'h57B8: data_out = 8'h1F;
                    16'h57B9: data_out = 8'h1E;
                    16'h57BA: data_out = 8'h1D;
                    16'h57BB: data_out = 8'h1C;
                    16'h57BC: data_out = 8'h1B;
                    16'h57BD: data_out = 8'h1A;
                    16'h57BE: data_out = 8'h19;
                    16'h57BF: data_out = 8'h18;
                    16'h57C0: data_out = 8'h17;
                    16'h57C1: data_out = 8'h16;
                    16'h57C2: data_out = 8'h15;
                    16'h57C3: data_out = 8'h14;
                    16'h57C4: data_out = 8'h13;
                    16'h57C5: data_out = 8'h12;
                    16'h57C6: data_out = 8'h11;
                    16'h57C7: data_out = 8'h10;
                    16'h57C8: data_out = 8'hF;
                    16'h57C9: data_out = 8'hE;
                    16'h57CA: data_out = 8'hD;
                    16'h57CB: data_out = 8'hC;
                    16'h57CC: data_out = 8'hB;
                    16'h57CD: data_out = 8'hA;
                    16'h57CE: data_out = 8'h9;
                    16'h57CF: data_out = 8'h8;
                    16'h57D0: data_out = 8'h7;
                    16'h57D1: data_out = 8'h6;
                    16'h57D2: data_out = 8'h5;
                    16'h57D3: data_out = 8'h4;
                    16'h57D4: data_out = 8'h3;
                    16'h57D5: data_out = 8'h2;
                    16'h57D6: data_out = 8'h1;
                    16'h57D7: data_out = 8'h0;
                    16'h57D8: data_out = 8'h81;
                    16'h57D9: data_out = 8'h82;
                    16'h57DA: data_out = 8'h83;
                    16'h57DB: data_out = 8'h84;
                    16'h57DC: data_out = 8'h85;
                    16'h57DD: data_out = 8'h86;
                    16'h57DE: data_out = 8'h87;
                    16'h57DF: data_out = 8'h88;
                    16'h57E0: data_out = 8'h89;
                    16'h57E1: data_out = 8'h8A;
                    16'h57E2: data_out = 8'h8B;
                    16'h57E3: data_out = 8'h8C;
                    16'h57E4: data_out = 8'h8D;
                    16'h57E5: data_out = 8'h8E;
                    16'h57E6: data_out = 8'h8F;
                    16'h57E7: data_out = 8'h90;
                    16'h57E8: data_out = 8'h91;
                    16'h57E9: data_out = 8'h92;
                    16'h57EA: data_out = 8'h93;
                    16'h57EB: data_out = 8'h94;
                    16'h57EC: data_out = 8'h95;
                    16'h57ED: data_out = 8'h96;
                    16'h57EE: data_out = 8'h97;
                    16'h57EF: data_out = 8'h98;
                    16'h57F0: data_out = 8'h99;
                    16'h57F1: data_out = 8'h9A;
                    16'h57F2: data_out = 8'h9B;
                    16'h57F3: data_out = 8'h9C;
                    16'h57F4: data_out = 8'h9D;
                    16'h57F5: data_out = 8'h9E;
                    16'h57F6: data_out = 8'h9F;
                    16'h57F7: data_out = 8'hA0;
                    16'h57F8: data_out = 8'hA1;
                    16'h57F9: data_out = 8'hA2;
                    16'h57FA: data_out = 8'hA3;
                    16'h57FB: data_out = 8'hA4;
                    16'h57FC: data_out = 8'hA5;
                    16'h57FD: data_out = 8'hA6;
                    16'h57FE: data_out = 8'hA7;
                    16'h57FF: data_out = 8'hA8;
                    16'h5800: data_out = 8'h58;
                    16'h5801: data_out = 8'h59;
                    16'h5802: data_out = 8'h5A;
                    16'h5803: data_out = 8'h5B;
                    16'h5804: data_out = 8'h5C;
                    16'h5805: data_out = 8'h5D;
                    16'h5806: data_out = 8'h5E;
                    16'h5807: data_out = 8'h5F;
                    16'h5808: data_out = 8'h60;
                    16'h5809: data_out = 8'h61;
                    16'h580A: data_out = 8'h62;
                    16'h580B: data_out = 8'h63;
                    16'h580C: data_out = 8'h64;
                    16'h580D: data_out = 8'h65;
                    16'h580E: data_out = 8'h66;
                    16'h580F: data_out = 8'h67;
                    16'h5810: data_out = 8'h68;
                    16'h5811: data_out = 8'h69;
                    16'h5812: data_out = 8'h6A;
                    16'h5813: data_out = 8'h6B;
                    16'h5814: data_out = 8'h6C;
                    16'h5815: data_out = 8'h6D;
                    16'h5816: data_out = 8'h6E;
                    16'h5817: data_out = 8'h6F;
                    16'h5818: data_out = 8'h70;
                    16'h5819: data_out = 8'h71;
                    16'h581A: data_out = 8'h72;
                    16'h581B: data_out = 8'h73;
                    16'h581C: data_out = 8'h74;
                    16'h581D: data_out = 8'h75;
                    16'h581E: data_out = 8'h76;
                    16'h581F: data_out = 8'h77;
                    16'h5820: data_out = 8'h78;
                    16'h5821: data_out = 8'h79;
                    16'h5822: data_out = 8'h7A;
                    16'h5823: data_out = 8'h7B;
                    16'h5824: data_out = 8'h7C;
                    16'h5825: data_out = 8'h7D;
                    16'h5826: data_out = 8'h7E;
                    16'h5827: data_out = 8'h7F;
                    16'h5828: data_out = 8'h80;
                    16'h5829: data_out = 8'h81;
                    16'h582A: data_out = 8'h82;
                    16'h582B: data_out = 8'h83;
                    16'h582C: data_out = 8'h84;
                    16'h582D: data_out = 8'h85;
                    16'h582E: data_out = 8'h86;
                    16'h582F: data_out = 8'h87;
                    16'h5830: data_out = 8'h88;
                    16'h5831: data_out = 8'h89;
                    16'h5832: data_out = 8'h8A;
                    16'h5833: data_out = 8'h8B;
                    16'h5834: data_out = 8'h8C;
                    16'h5835: data_out = 8'h8D;
                    16'h5836: data_out = 8'h8E;
                    16'h5837: data_out = 8'h8F;
                    16'h5838: data_out = 8'h90;
                    16'h5839: data_out = 8'h91;
                    16'h583A: data_out = 8'h92;
                    16'h583B: data_out = 8'h93;
                    16'h583C: data_out = 8'h94;
                    16'h583D: data_out = 8'h95;
                    16'h583E: data_out = 8'h96;
                    16'h583F: data_out = 8'h97;
                    16'h5840: data_out = 8'h98;
                    16'h5841: data_out = 8'h99;
                    16'h5842: data_out = 8'h9A;
                    16'h5843: data_out = 8'h9B;
                    16'h5844: data_out = 8'h9C;
                    16'h5845: data_out = 8'h9D;
                    16'h5846: data_out = 8'h9E;
                    16'h5847: data_out = 8'h9F;
                    16'h5848: data_out = 8'hA0;
                    16'h5849: data_out = 8'hA1;
                    16'h584A: data_out = 8'hA2;
                    16'h584B: data_out = 8'hA3;
                    16'h584C: data_out = 8'hA4;
                    16'h584D: data_out = 8'hA5;
                    16'h584E: data_out = 8'hA6;
                    16'h584F: data_out = 8'hA7;
                    16'h5850: data_out = 8'hA8;
                    16'h5851: data_out = 8'hA9;
                    16'h5852: data_out = 8'hAA;
                    16'h5853: data_out = 8'hAB;
                    16'h5854: data_out = 8'hAC;
                    16'h5855: data_out = 8'hAD;
                    16'h5856: data_out = 8'hAE;
                    16'h5857: data_out = 8'hAF;
                    16'h5858: data_out = 8'hB0;
                    16'h5859: data_out = 8'hB1;
                    16'h585A: data_out = 8'hB2;
                    16'h585B: data_out = 8'hB3;
                    16'h585C: data_out = 8'hB4;
                    16'h585D: data_out = 8'hB5;
                    16'h585E: data_out = 8'hB6;
                    16'h585F: data_out = 8'hB7;
                    16'h5860: data_out = 8'hB8;
                    16'h5861: data_out = 8'hB9;
                    16'h5862: data_out = 8'hBA;
                    16'h5863: data_out = 8'hBB;
                    16'h5864: data_out = 8'hBC;
                    16'h5865: data_out = 8'hBD;
                    16'h5866: data_out = 8'hBE;
                    16'h5867: data_out = 8'hBF;
                    16'h5868: data_out = 8'hC0;
                    16'h5869: data_out = 8'hC1;
                    16'h586A: data_out = 8'hC2;
                    16'h586B: data_out = 8'hC3;
                    16'h586C: data_out = 8'hC4;
                    16'h586D: data_out = 8'hC5;
                    16'h586E: data_out = 8'hC6;
                    16'h586F: data_out = 8'hC7;
                    16'h5870: data_out = 8'hC8;
                    16'h5871: data_out = 8'hC9;
                    16'h5872: data_out = 8'hCA;
                    16'h5873: data_out = 8'hCB;
                    16'h5874: data_out = 8'hCC;
                    16'h5875: data_out = 8'hCD;
                    16'h5876: data_out = 8'hCE;
                    16'h5877: data_out = 8'hCF;
                    16'h5878: data_out = 8'hD0;
                    16'h5879: data_out = 8'hD1;
                    16'h587A: data_out = 8'hD2;
                    16'h587B: data_out = 8'hD3;
                    16'h587C: data_out = 8'hD4;
                    16'h587D: data_out = 8'hD5;
                    16'h587E: data_out = 8'hD6;
                    16'h587F: data_out = 8'hD7;
                    16'h5880: data_out = 8'h58;
                    16'h5881: data_out = 8'h57;
                    16'h5882: data_out = 8'h56;
                    16'h5883: data_out = 8'h55;
                    16'h5884: data_out = 8'h54;
                    16'h5885: data_out = 8'h53;
                    16'h5886: data_out = 8'h52;
                    16'h5887: data_out = 8'h51;
                    16'h5888: data_out = 8'h50;
                    16'h5889: data_out = 8'h4F;
                    16'h588A: data_out = 8'h4E;
                    16'h588B: data_out = 8'h4D;
                    16'h588C: data_out = 8'h4C;
                    16'h588D: data_out = 8'h4B;
                    16'h588E: data_out = 8'h4A;
                    16'h588F: data_out = 8'h49;
                    16'h5890: data_out = 8'h48;
                    16'h5891: data_out = 8'h47;
                    16'h5892: data_out = 8'h46;
                    16'h5893: data_out = 8'h45;
                    16'h5894: data_out = 8'h44;
                    16'h5895: data_out = 8'h43;
                    16'h5896: data_out = 8'h42;
                    16'h5897: data_out = 8'h41;
                    16'h5898: data_out = 8'h40;
                    16'h5899: data_out = 8'h3F;
                    16'h589A: data_out = 8'h3E;
                    16'h589B: data_out = 8'h3D;
                    16'h589C: data_out = 8'h3C;
                    16'h589D: data_out = 8'h3B;
                    16'h589E: data_out = 8'h3A;
                    16'h589F: data_out = 8'h39;
                    16'h58A0: data_out = 8'h38;
                    16'h58A1: data_out = 8'h37;
                    16'h58A2: data_out = 8'h36;
                    16'h58A3: data_out = 8'h35;
                    16'h58A4: data_out = 8'h34;
                    16'h58A5: data_out = 8'h33;
                    16'h58A6: data_out = 8'h32;
                    16'h58A7: data_out = 8'h31;
                    16'h58A8: data_out = 8'h30;
                    16'h58A9: data_out = 8'h2F;
                    16'h58AA: data_out = 8'h2E;
                    16'h58AB: data_out = 8'h2D;
                    16'h58AC: data_out = 8'h2C;
                    16'h58AD: data_out = 8'h2B;
                    16'h58AE: data_out = 8'h2A;
                    16'h58AF: data_out = 8'h29;
                    16'h58B0: data_out = 8'h28;
                    16'h58B1: data_out = 8'h27;
                    16'h58B2: data_out = 8'h26;
                    16'h58B3: data_out = 8'h25;
                    16'h58B4: data_out = 8'h24;
                    16'h58B5: data_out = 8'h23;
                    16'h58B6: data_out = 8'h22;
                    16'h58B7: data_out = 8'h21;
                    16'h58B8: data_out = 8'h20;
                    16'h58B9: data_out = 8'h1F;
                    16'h58BA: data_out = 8'h1E;
                    16'h58BB: data_out = 8'h1D;
                    16'h58BC: data_out = 8'h1C;
                    16'h58BD: data_out = 8'h1B;
                    16'h58BE: data_out = 8'h1A;
                    16'h58BF: data_out = 8'h19;
                    16'h58C0: data_out = 8'h18;
                    16'h58C1: data_out = 8'h17;
                    16'h58C2: data_out = 8'h16;
                    16'h58C3: data_out = 8'h15;
                    16'h58C4: data_out = 8'h14;
                    16'h58C5: data_out = 8'h13;
                    16'h58C6: data_out = 8'h12;
                    16'h58C7: data_out = 8'h11;
                    16'h58C8: data_out = 8'h10;
                    16'h58C9: data_out = 8'hF;
                    16'h58CA: data_out = 8'hE;
                    16'h58CB: data_out = 8'hD;
                    16'h58CC: data_out = 8'hC;
                    16'h58CD: data_out = 8'hB;
                    16'h58CE: data_out = 8'hA;
                    16'h58CF: data_out = 8'h9;
                    16'h58D0: data_out = 8'h8;
                    16'h58D1: data_out = 8'h7;
                    16'h58D2: data_out = 8'h6;
                    16'h58D3: data_out = 8'h5;
                    16'h58D4: data_out = 8'h4;
                    16'h58D5: data_out = 8'h3;
                    16'h58D6: data_out = 8'h2;
                    16'h58D7: data_out = 8'h1;
                    16'h58D8: data_out = 8'h0;
                    16'h58D9: data_out = 8'h81;
                    16'h58DA: data_out = 8'h82;
                    16'h58DB: data_out = 8'h83;
                    16'h58DC: data_out = 8'h84;
                    16'h58DD: data_out = 8'h85;
                    16'h58DE: data_out = 8'h86;
                    16'h58DF: data_out = 8'h87;
                    16'h58E0: data_out = 8'h88;
                    16'h58E1: data_out = 8'h89;
                    16'h58E2: data_out = 8'h8A;
                    16'h58E3: data_out = 8'h8B;
                    16'h58E4: data_out = 8'h8C;
                    16'h58E5: data_out = 8'h8D;
                    16'h58E6: data_out = 8'h8E;
                    16'h58E7: data_out = 8'h8F;
                    16'h58E8: data_out = 8'h90;
                    16'h58E9: data_out = 8'h91;
                    16'h58EA: data_out = 8'h92;
                    16'h58EB: data_out = 8'h93;
                    16'h58EC: data_out = 8'h94;
                    16'h58ED: data_out = 8'h95;
                    16'h58EE: data_out = 8'h96;
                    16'h58EF: data_out = 8'h97;
                    16'h58F0: data_out = 8'h98;
                    16'h58F1: data_out = 8'h99;
                    16'h58F2: data_out = 8'h9A;
                    16'h58F3: data_out = 8'h9B;
                    16'h58F4: data_out = 8'h9C;
                    16'h58F5: data_out = 8'h9D;
                    16'h58F6: data_out = 8'h9E;
                    16'h58F7: data_out = 8'h9F;
                    16'h58F8: data_out = 8'hA0;
                    16'h58F9: data_out = 8'hA1;
                    16'h58FA: data_out = 8'hA2;
                    16'h58FB: data_out = 8'hA3;
                    16'h58FC: data_out = 8'hA4;
                    16'h58FD: data_out = 8'hA5;
                    16'h58FE: data_out = 8'hA6;
                    16'h58FF: data_out = 8'hA7;
                    16'h5900: data_out = 8'h59;
                    16'h5901: data_out = 8'h5A;
                    16'h5902: data_out = 8'h5B;
                    16'h5903: data_out = 8'h5C;
                    16'h5904: data_out = 8'h5D;
                    16'h5905: data_out = 8'h5E;
                    16'h5906: data_out = 8'h5F;
                    16'h5907: data_out = 8'h60;
                    16'h5908: data_out = 8'h61;
                    16'h5909: data_out = 8'h62;
                    16'h590A: data_out = 8'h63;
                    16'h590B: data_out = 8'h64;
                    16'h590C: data_out = 8'h65;
                    16'h590D: data_out = 8'h66;
                    16'h590E: data_out = 8'h67;
                    16'h590F: data_out = 8'h68;
                    16'h5910: data_out = 8'h69;
                    16'h5911: data_out = 8'h6A;
                    16'h5912: data_out = 8'h6B;
                    16'h5913: data_out = 8'h6C;
                    16'h5914: data_out = 8'h6D;
                    16'h5915: data_out = 8'h6E;
                    16'h5916: data_out = 8'h6F;
                    16'h5917: data_out = 8'h70;
                    16'h5918: data_out = 8'h71;
                    16'h5919: data_out = 8'h72;
                    16'h591A: data_out = 8'h73;
                    16'h591B: data_out = 8'h74;
                    16'h591C: data_out = 8'h75;
                    16'h591D: data_out = 8'h76;
                    16'h591E: data_out = 8'h77;
                    16'h591F: data_out = 8'h78;
                    16'h5920: data_out = 8'h79;
                    16'h5921: data_out = 8'h7A;
                    16'h5922: data_out = 8'h7B;
                    16'h5923: data_out = 8'h7C;
                    16'h5924: data_out = 8'h7D;
                    16'h5925: data_out = 8'h7E;
                    16'h5926: data_out = 8'h7F;
                    16'h5927: data_out = 8'h80;
                    16'h5928: data_out = 8'h81;
                    16'h5929: data_out = 8'h82;
                    16'h592A: data_out = 8'h83;
                    16'h592B: data_out = 8'h84;
                    16'h592C: data_out = 8'h85;
                    16'h592D: data_out = 8'h86;
                    16'h592E: data_out = 8'h87;
                    16'h592F: data_out = 8'h88;
                    16'h5930: data_out = 8'h89;
                    16'h5931: data_out = 8'h8A;
                    16'h5932: data_out = 8'h8B;
                    16'h5933: data_out = 8'h8C;
                    16'h5934: data_out = 8'h8D;
                    16'h5935: data_out = 8'h8E;
                    16'h5936: data_out = 8'h8F;
                    16'h5937: data_out = 8'h90;
                    16'h5938: data_out = 8'h91;
                    16'h5939: data_out = 8'h92;
                    16'h593A: data_out = 8'h93;
                    16'h593B: data_out = 8'h94;
                    16'h593C: data_out = 8'h95;
                    16'h593D: data_out = 8'h96;
                    16'h593E: data_out = 8'h97;
                    16'h593F: data_out = 8'h98;
                    16'h5940: data_out = 8'h99;
                    16'h5941: data_out = 8'h9A;
                    16'h5942: data_out = 8'h9B;
                    16'h5943: data_out = 8'h9C;
                    16'h5944: data_out = 8'h9D;
                    16'h5945: data_out = 8'h9E;
                    16'h5946: data_out = 8'h9F;
                    16'h5947: data_out = 8'hA0;
                    16'h5948: data_out = 8'hA1;
                    16'h5949: data_out = 8'hA2;
                    16'h594A: data_out = 8'hA3;
                    16'h594B: data_out = 8'hA4;
                    16'h594C: data_out = 8'hA5;
                    16'h594D: data_out = 8'hA6;
                    16'h594E: data_out = 8'hA7;
                    16'h594F: data_out = 8'hA8;
                    16'h5950: data_out = 8'hA9;
                    16'h5951: data_out = 8'hAA;
                    16'h5952: data_out = 8'hAB;
                    16'h5953: data_out = 8'hAC;
                    16'h5954: data_out = 8'hAD;
                    16'h5955: data_out = 8'hAE;
                    16'h5956: data_out = 8'hAF;
                    16'h5957: data_out = 8'hB0;
                    16'h5958: data_out = 8'hB1;
                    16'h5959: data_out = 8'hB2;
                    16'h595A: data_out = 8'hB3;
                    16'h595B: data_out = 8'hB4;
                    16'h595C: data_out = 8'hB5;
                    16'h595D: data_out = 8'hB6;
                    16'h595E: data_out = 8'hB7;
                    16'h595F: data_out = 8'hB8;
                    16'h5960: data_out = 8'hB9;
                    16'h5961: data_out = 8'hBA;
                    16'h5962: data_out = 8'hBB;
                    16'h5963: data_out = 8'hBC;
                    16'h5964: data_out = 8'hBD;
                    16'h5965: data_out = 8'hBE;
                    16'h5966: data_out = 8'hBF;
                    16'h5967: data_out = 8'hC0;
                    16'h5968: data_out = 8'hC1;
                    16'h5969: data_out = 8'hC2;
                    16'h596A: data_out = 8'hC3;
                    16'h596B: data_out = 8'hC4;
                    16'h596C: data_out = 8'hC5;
                    16'h596D: data_out = 8'hC6;
                    16'h596E: data_out = 8'hC7;
                    16'h596F: data_out = 8'hC8;
                    16'h5970: data_out = 8'hC9;
                    16'h5971: data_out = 8'hCA;
                    16'h5972: data_out = 8'hCB;
                    16'h5973: data_out = 8'hCC;
                    16'h5974: data_out = 8'hCD;
                    16'h5975: data_out = 8'hCE;
                    16'h5976: data_out = 8'hCF;
                    16'h5977: data_out = 8'hD0;
                    16'h5978: data_out = 8'hD1;
                    16'h5979: data_out = 8'hD2;
                    16'h597A: data_out = 8'hD3;
                    16'h597B: data_out = 8'hD4;
                    16'h597C: data_out = 8'hD5;
                    16'h597D: data_out = 8'hD6;
                    16'h597E: data_out = 8'hD7;
                    16'h597F: data_out = 8'hD8;
                    16'h5980: data_out = 8'h59;
                    16'h5981: data_out = 8'h58;
                    16'h5982: data_out = 8'h57;
                    16'h5983: data_out = 8'h56;
                    16'h5984: data_out = 8'h55;
                    16'h5985: data_out = 8'h54;
                    16'h5986: data_out = 8'h53;
                    16'h5987: data_out = 8'h52;
                    16'h5988: data_out = 8'h51;
                    16'h5989: data_out = 8'h50;
                    16'h598A: data_out = 8'h4F;
                    16'h598B: data_out = 8'h4E;
                    16'h598C: data_out = 8'h4D;
                    16'h598D: data_out = 8'h4C;
                    16'h598E: data_out = 8'h4B;
                    16'h598F: data_out = 8'h4A;
                    16'h5990: data_out = 8'h49;
                    16'h5991: data_out = 8'h48;
                    16'h5992: data_out = 8'h47;
                    16'h5993: data_out = 8'h46;
                    16'h5994: data_out = 8'h45;
                    16'h5995: data_out = 8'h44;
                    16'h5996: data_out = 8'h43;
                    16'h5997: data_out = 8'h42;
                    16'h5998: data_out = 8'h41;
                    16'h5999: data_out = 8'h40;
                    16'h599A: data_out = 8'h3F;
                    16'h599B: data_out = 8'h3E;
                    16'h599C: data_out = 8'h3D;
                    16'h599D: data_out = 8'h3C;
                    16'h599E: data_out = 8'h3B;
                    16'h599F: data_out = 8'h3A;
                    16'h59A0: data_out = 8'h39;
                    16'h59A1: data_out = 8'h38;
                    16'h59A2: data_out = 8'h37;
                    16'h59A3: data_out = 8'h36;
                    16'h59A4: data_out = 8'h35;
                    16'h59A5: data_out = 8'h34;
                    16'h59A6: data_out = 8'h33;
                    16'h59A7: data_out = 8'h32;
                    16'h59A8: data_out = 8'h31;
                    16'h59A9: data_out = 8'h30;
                    16'h59AA: data_out = 8'h2F;
                    16'h59AB: data_out = 8'h2E;
                    16'h59AC: data_out = 8'h2D;
                    16'h59AD: data_out = 8'h2C;
                    16'h59AE: data_out = 8'h2B;
                    16'h59AF: data_out = 8'h2A;
                    16'h59B0: data_out = 8'h29;
                    16'h59B1: data_out = 8'h28;
                    16'h59B2: data_out = 8'h27;
                    16'h59B3: data_out = 8'h26;
                    16'h59B4: data_out = 8'h25;
                    16'h59B5: data_out = 8'h24;
                    16'h59B6: data_out = 8'h23;
                    16'h59B7: data_out = 8'h22;
                    16'h59B8: data_out = 8'h21;
                    16'h59B9: data_out = 8'h20;
                    16'h59BA: data_out = 8'h1F;
                    16'h59BB: data_out = 8'h1E;
                    16'h59BC: data_out = 8'h1D;
                    16'h59BD: data_out = 8'h1C;
                    16'h59BE: data_out = 8'h1B;
                    16'h59BF: data_out = 8'h1A;
                    16'h59C0: data_out = 8'h19;
                    16'h59C1: data_out = 8'h18;
                    16'h59C2: data_out = 8'h17;
                    16'h59C3: data_out = 8'h16;
                    16'h59C4: data_out = 8'h15;
                    16'h59C5: data_out = 8'h14;
                    16'h59C6: data_out = 8'h13;
                    16'h59C7: data_out = 8'h12;
                    16'h59C8: data_out = 8'h11;
                    16'h59C9: data_out = 8'h10;
                    16'h59CA: data_out = 8'hF;
                    16'h59CB: data_out = 8'hE;
                    16'h59CC: data_out = 8'hD;
                    16'h59CD: data_out = 8'hC;
                    16'h59CE: data_out = 8'hB;
                    16'h59CF: data_out = 8'hA;
                    16'h59D0: data_out = 8'h9;
                    16'h59D1: data_out = 8'h8;
                    16'h59D2: data_out = 8'h7;
                    16'h59D3: data_out = 8'h6;
                    16'h59D4: data_out = 8'h5;
                    16'h59D5: data_out = 8'h4;
                    16'h59D6: data_out = 8'h3;
                    16'h59D7: data_out = 8'h2;
                    16'h59D8: data_out = 8'h1;
                    16'h59D9: data_out = 8'h0;
                    16'h59DA: data_out = 8'h81;
                    16'h59DB: data_out = 8'h82;
                    16'h59DC: data_out = 8'h83;
                    16'h59DD: data_out = 8'h84;
                    16'h59DE: data_out = 8'h85;
                    16'h59DF: data_out = 8'h86;
                    16'h59E0: data_out = 8'h87;
                    16'h59E1: data_out = 8'h88;
                    16'h59E2: data_out = 8'h89;
                    16'h59E3: data_out = 8'h8A;
                    16'h59E4: data_out = 8'h8B;
                    16'h59E5: data_out = 8'h8C;
                    16'h59E6: data_out = 8'h8D;
                    16'h59E7: data_out = 8'h8E;
                    16'h59E8: data_out = 8'h8F;
                    16'h59E9: data_out = 8'h90;
                    16'h59EA: data_out = 8'h91;
                    16'h59EB: data_out = 8'h92;
                    16'h59EC: data_out = 8'h93;
                    16'h59ED: data_out = 8'h94;
                    16'h59EE: data_out = 8'h95;
                    16'h59EF: data_out = 8'h96;
                    16'h59F0: data_out = 8'h97;
                    16'h59F1: data_out = 8'h98;
                    16'h59F2: data_out = 8'h99;
                    16'h59F3: data_out = 8'h9A;
                    16'h59F4: data_out = 8'h9B;
                    16'h59F5: data_out = 8'h9C;
                    16'h59F6: data_out = 8'h9D;
                    16'h59F7: data_out = 8'h9E;
                    16'h59F8: data_out = 8'h9F;
                    16'h59F9: data_out = 8'hA0;
                    16'h59FA: data_out = 8'hA1;
                    16'h59FB: data_out = 8'hA2;
                    16'h59FC: data_out = 8'hA3;
                    16'h59FD: data_out = 8'hA4;
                    16'h59FE: data_out = 8'hA5;
                    16'h59FF: data_out = 8'hA6;
                    16'h5A00: data_out = 8'h5A;
                    16'h5A01: data_out = 8'h5B;
                    16'h5A02: data_out = 8'h5C;
                    16'h5A03: data_out = 8'h5D;
                    16'h5A04: data_out = 8'h5E;
                    16'h5A05: data_out = 8'h5F;
                    16'h5A06: data_out = 8'h60;
                    16'h5A07: data_out = 8'h61;
                    16'h5A08: data_out = 8'h62;
                    16'h5A09: data_out = 8'h63;
                    16'h5A0A: data_out = 8'h64;
                    16'h5A0B: data_out = 8'h65;
                    16'h5A0C: data_out = 8'h66;
                    16'h5A0D: data_out = 8'h67;
                    16'h5A0E: data_out = 8'h68;
                    16'h5A0F: data_out = 8'h69;
                    16'h5A10: data_out = 8'h6A;
                    16'h5A11: data_out = 8'h6B;
                    16'h5A12: data_out = 8'h6C;
                    16'h5A13: data_out = 8'h6D;
                    16'h5A14: data_out = 8'h6E;
                    16'h5A15: data_out = 8'h6F;
                    16'h5A16: data_out = 8'h70;
                    16'h5A17: data_out = 8'h71;
                    16'h5A18: data_out = 8'h72;
                    16'h5A19: data_out = 8'h73;
                    16'h5A1A: data_out = 8'h74;
                    16'h5A1B: data_out = 8'h75;
                    16'h5A1C: data_out = 8'h76;
                    16'h5A1D: data_out = 8'h77;
                    16'h5A1E: data_out = 8'h78;
                    16'h5A1F: data_out = 8'h79;
                    16'h5A20: data_out = 8'h7A;
                    16'h5A21: data_out = 8'h7B;
                    16'h5A22: data_out = 8'h7C;
                    16'h5A23: data_out = 8'h7D;
                    16'h5A24: data_out = 8'h7E;
                    16'h5A25: data_out = 8'h7F;
                    16'h5A26: data_out = 8'h80;
                    16'h5A27: data_out = 8'h81;
                    16'h5A28: data_out = 8'h82;
                    16'h5A29: data_out = 8'h83;
                    16'h5A2A: data_out = 8'h84;
                    16'h5A2B: data_out = 8'h85;
                    16'h5A2C: data_out = 8'h86;
                    16'h5A2D: data_out = 8'h87;
                    16'h5A2E: data_out = 8'h88;
                    16'h5A2F: data_out = 8'h89;
                    16'h5A30: data_out = 8'h8A;
                    16'h5A31: data_out = 8'h8B;
                    16'h5A32: data_out = 8'h8C;
                    16'h5A33: data_out = 8'h8D;
                    16'h5A34: data_out = 8'h8E;
                    16'h5A35: data_out = 8'h8F;
                    16'h5A36: data_out = 8'h90;
                    16'h5A37: data_out = 8'h91;
                    16'h5A38: data_out = 8'h92;
                    16'h5A39: data_out = 8'h93;
                    16'h5A3A: data_out = 8'h94;
                    16'h5A3B: data_out = 8'h95;
                    16'h5A3C: data_out = 8'h96;
                    16'h5A3D: data_out = 8'h97;
                    16'h5A3E: data_out = 8'h98;
                    16'h5A3F: data_out = 8'h99;
                    16'h5A40: data_out = 8'h9A;
                    16'h5A41: data_out = 8'h9B;
                    16'h5A42: data_out = 8'h9C;
                    16'h5A43: data_out = 8'h9D;
                    16'h5A44: data_out = 8'h9E;
                    16'h5A45: data_out = 8'h9F;
                    16'h5A46: data_out = 8'hA0;
                    16'h5A47: data_out = 8'hA1;
                    16'h5A48: data_out = 8'hA2;
                    16'h5A49: data_out = 8'hA3;
                    16'h5A4A: data_out = 8'hA4;
                    16'h5A4B: data_out = 8'hA5;
                    16'h5A4C: data_out = 8'hA6;
                    16'h5A4D: data_out = 8'hA7;
                    16'h5A4E: data_out = 8'hA8;
                    16'h5A4F: data_out = 8'hA9;
                    16'h5A50: data_out = 8'hAA;
                    16'h5A51: data_out = 8'hAB;
                    16'h5A52: data_out = 8'hAC;
                    16'h5A53: data_out = 8'hAD;
                    16'h5A54: data_out = 8'hAE;
                    16'h5A55: data_out = 8'hAF;
                    16'h5A56: data_out = 8'hB0;
                    16'h5A57: data_out = 8'hB1;
                    16'h5A58: data_out = 8'hB2;
                    16'h5A59: data_out = 8'hB3;
                    16'h5A5A: data_out = 8'hB4;
                    16'h5A5B: data_out = 8'hB5;
                    16'h5A5C: data_out = 8'hB6;
                    16'h5A5D: data_out = 8'hB7;
                    16'h5A5E: data_out = 8'hB8;
                    16'h5A5F: data_out = 8'hB9;
                    16'h5A60: data_out = 8'hBA;
                    16'h5A61: data_out = 8'hBB;
                    16'h5A62: data_out = 8'hBC;
                    16'h5A63: data_out = 8'hBD;
                    16'h5A64: data_out = 8'hBE;
                    16'h5A65: data_out = 8'hBF;
                    16'h5A66: data_out = 8'hC0;
                    16'h5A67: data_out = 8'hC1;
                    16'h5A68: data_out = 8'hC2;
                    16'h5A69: data_out = 8'hC3;
                    16'h5A6A: data_out = 8'hC4;
                    16'h5A6B: data_out = 8'hC5;
                    16'h5A6C: data_out = 8'hC6;
                    16'h5A6D: data_out = 8'hC7;
                    16'h5A6E: data_out = 8'hC8;
                    16'h5A6F: data_out = 8'hC9;
                    16'h5A70: data_out = 8'hCA;
                    16'h5A71: data_out = 8'hCB;
                    16'h5A72: data_out = 8'hCC;
                    16'h5A73: data_out = 8'hCD;
                    16'h5A74: data_out = 8'hCE;
                    16'h5A75: data_out = 8'hCF;
                    16'h5A76: data_out = 8'hD0;
                    16'h5A77: data_out = 8'hD1;
                    16'h5A78: data_out = 8'hD2;
                    16'h5A79: data_out = 8'hD3;
                    16'h5A7A: data_out = 8'hD4;
                    16'h5A7B: data_out = 8'hD5;
                    16'h5A7C: data_out = 8'hD6;
                    16'h5A7D: data_out = 8'hD7;
                    16'h5A7E: data_out = 8'hD8;
                    16'h5A7F: data_out = 8'hD9;
                    16'h5A80: data_out = 8'h5A;
                    16'h5A81: data_out = 8'h59;
                    16'h5A82: data_out = 8'h58;
                    16'h5A83: data_out = 8'h57;
                    16'h5A84: data_out = 8'h56;
                    16'h5A85: data_out = 8'h55;
                    16'h5A86: data_out = 8'h54;
                    16'h5A87: data_out = 8'h53;
                    16'h5A88: data_out = 8'h52;
                    16'h5A89: data_out = 8'h51;
                    16'h5A8A: data_out = 8'h50;
                    16'h5A8B: data_out = 8'h4F;
                    16'h5A8C: data_out = 8'h4E;
                    16'h5A8D: data_out = 8'h4D;
                    16'h5A8E: data_out = 8'h4C;
                    16'h5A8F: data_out = 8'h4B;
                    16'h5A90: data_out = 8'h4A;
                    16'h5A91: data_out = 8'h49;
                    16'h5A92: data_out = 8'h48;
                    16'h5A93: data_out = 8'h47;
                    16'h5A94: data_out = 8'h46;
                    16'h5A95: data_out = 8'h45;
                    16'h5A96: data_out = 8'h44;
                    16'h5A97: data_out = 8'h43;
                    16'h5A98: data_out = 8'h42;
                    16'h5A99: data_out = 8'h41;
                    16'h5A9A: data_out = 8'h40;
                    16'h5A9B: data_out = 8'h3F;
                    16'h5A9C: data_out = 8'h3E;
                    16'h5A9D: data_out = 8'h3D;
                    16'h5A9E: data_out = 8'h3C;
                    16'h5A9F: data_out = 8'h3B;
                    16'h5AA0: data_out = 8'h3A;
                    16'h5AA1: data_out = 8'h39;
                    16'h5AA2: data_out = 8'h38;
                    16'h5AA3: data_out = 8'h37;
                    16'h5AA4: data_out = 8'h36;
                    16'h5AA5: data_out = 8'h35;
                    16'h5AA6: data_out = 8'h34;
                    16'h5AA7: data_out = 8'h33;
                    16'h5AA8: data_out = 8'h32;
                    16'h5AA9: data_out = 8'h31;
                    16'h5AAA: data_out = 8'h30;
                    16'h5AAB: data_out = 8'h2F;
                    16'h5AAC: data_out = 8'h2E;
                    16'h5AAD: data_out = 8'h2D;
                    16'h5AAE: data_out = 8'h2C;
                    16'h5AAF: data_out = 8'h2B;
                    16'h5AB0: data_out = 8'h2A;
                    16'h5AB1: data_out = 8'h29;
                    16'h5AB2: data_out = 8'h28;
                    16'h5AB3: data_out = 8'h27;
                    16'h5AB4: data_out = 8'h26;
                    16'h5AB5: data_out = 8'h25;
                    16'h5AB6: data_out = 8'h24;
                    16'h5AB7: data_out = 8'h23;
                    16'h5AB8: data_out = 8'h22;
                    16'h5AB9: data_out = 8'h21;
                    16'h5ABA: data_out = 8'h20;
                    16'h5ABB: data_out = 8'h1F;
                    16'h5ABC: data_out = 8'h1E;
                    16'h5ABD: data_out = 8'h1D;
                    16'h5ABE: data_out = 8'h1C;
                    16'h5ABF: data_out = 8'h1B;
                    16'h5AC0: data_out = 8'h1A;
                    16'h5AC1: data_out = 8'h19;
                    16'h5AC2: data_out = 8'h18;
                    16'h5AC3: data_out = 8'h17;
                    16'h5AC4: data_out = 8'h16;
                    16'h5AC5: data_out = 8'h15;
                    16'h5AC6: data_out = 8'h14;
                    16'h5AC7: data_out = 8'h13;
                    16'h5AC8: data_out = 8'h12;
                    16'h5AC9: data_out = 8'h11;
                    16'h5ACA: data_out = 8'h10;
                    16'h5ACB: data_out = 8'hF;
                    16'h5ACC: data_out = 8'hE;
                    16'h5ACD: data_out = 8'hD;
                    16'h5ACE: data_out = 8'hC;
                    16'h5ACF: data_out = 8'hB;
                    16'h5AD0: data_out = 8'hA;
                    16'h5AD1: data_out = 8'h9;
                    16'h5AD2: data_out = 8'h8;
                    16'h5AD3: data_out = 8'h7;
                    16'h5AD4: data_out = 8'h6;
                    16'h5AD5: data_out = 8'h5;
                    16'h5AD6: data_out = 8'h4;
                    16'h5AD7: data_out = 8'h3;
                    16'h5AD8: data_out = 8'h2;
                    16'h5AD9: data_out = 8'h1;
                    16'h5ADA: data_out = 8'h0;
                    16'h5ADB: data_out = 8'h81;
                    16'h5ADC: data_out = 8'h82;
                    16'h5ADD: data_out = 8'h83;
                    16'h5ADE: data_out = 8'h84;
                    16'h5ADF: data_out = 8'h85;
                    16'h5AE0: data_out = 8'h86;
                    16'h5AE1: data_out = 8'h87;
                    16'h5AE2: data_out = 8'h88;
                    16'h5AE3: data_out = 8'h89;
                    16'h5AE4: data_out = 8'h8A;
                    16'h5AE5: data_out = 8'h8B;
                    16'h5AE6: data_out = 8'h8C;
                    16'h5AE7: data_out = 8'h8D;
                    16'h5AE8: data_out = 8'h8E;
                    16'h5AE9: data_out = 8'h8F;
                    16'h5AEA: data_out = 8'h90;
                    16'h5AEB: data_out = 8'h91;
                    16'h5AEC: data_out = 8'h92;
                    16'h5AED: data_out = 8'h93;
                    16'h5AEE: data_out = 8'h94;
                    16'h5AEF: data_out = 8'h95;
                    16'h5AF0: data_out = 8'h96;
                    16'h5AF1: data_out = 8'h97;
                    16'h5AF2: data_out = 8'h98;
                    16'h5AF3: data_out = 8'h99;
                    16'h5AF4: data_out = 8'h9A;
                    16'h5AF5: data_out = 8'h9B;
                    16'h5AF6: data_out = 8'h9C;
                    16'h5AF7: data_out = 8'h9D;
                    16'h5AF8: data_out = 8'h9E;
                    16'h5AF9: data_out = 8'h9F;
                    16'h5AFA: data_out = 8'hA0;
                    16'h5AFB: data_out = 8'hA1;
                    16'h5AFC: data_out = 8'hA2;
                    16'h5AFD: data_out = 8'hA3;
                    16'h5AFE: data_out = 8'hA4;
                    16'h5AFF: data_out = 8'hA5;
                    16'h5B00: data_out = 8'h5B;
                    16'h5B01: data_out = 8'h5C;
                    16'h5B02: data_out = 8'h5D;
                    16'h5B03: data_out = 8'h5E;
                    16'h5B04: data_out = 8'h5F;
                    16'h5B05: data_out = 8'h60;
                    16'h5B06: data_out = 8'h61;
                    16'h5B07: data_out = 8'h62;
                    16'h5B08: data_out = 8'h63;
                    16'h5B09: data_out = 8'h64;
                    16'h5B0A: data_out = 8'h65;
                    16'h5B0B: data_out = 8'h66;
                    16'h5B0C: data_out = 8'h67;
                    16'h5B0D: data_out = 8'h68;
                    16'h5B0E: data_out = 8'h69;
                    16'h5B0F: data_out = 8'h6A;
                    16'h5B10: data_out = 8'h6B;
                    16'h5B11: data_out = 8'h6C;
                    16'h5B12: data_out = 8'h6D;
                    16'h5B13: data_out = 8'h6E;
                    16'h5B14: data_out = 8'h6F;
                    16'h5B15: data_out = 8'h70;
                    16'h5B16: data_out = 8'h71;
                    16'h5B17: data_out = 8'h72;
                    16'h5B18: data_out = 8'h73;
                    16'h5B19: data_out = 8'h74;
                    16'h5B1A: data_out = 8'h75;
                    16'h5B1B: data_out = 8'h76;
                    16'h5B1C: data_out = 8'h77;
                    16'h5B1D: data_out = 8'h78;
                    16'h5B1E: data_out = 8'h79;
                    16'h5B1F: data_out = 8'h7A;
                    16'h5B20: data_out = 8'h7B;
                    16'h5B21: data_out = 8'h7C;
                    16'h5B22: data_out = 8'h7D;
                    16'h5B23: data_out = 8'h7E;
                    16'h5B24: data_out = 8'h7F;
                    16'h5B25: data_out = 8'h80;
                    16'h5B26: data_out = 8'h81;
                    16'h5B27: data_out = 8'h82;
                    16'h5B28: data_out = 8'h83;
                    16'h5B29: data_out = 8'h84;
                    16'h5B2A: data_out = 8'h85;
                    16'h5B2B: data_out = 8'h86;
                    16'h5B2C: data_out = 8'h87;
                    16'h5B2D: data_out = 8'h88;
                    16'h5B2E: data_out = 8'h89;
                    16'h5B2F: data_out = 8'h8A;
                    16'h5B30: data_out = 8'h8B;
                    16'h5B31: data_out = 8'h8C;
                    16'h5B32: data_out = 8'h8D;
                    16'h5B33: data_out = 8'h8E;
                    16'h5B34: data_out = 8'h8F;
                    16'h5B35: data_out = 8'h90;
                    16'h5B36: data_out = 8'h91;
                    16'h5B37: data_out = 8'h92;
                    16'h5B38: data_out = 8'h93;
                    16'h5B39: data_out = 8'h94;
                    16'h5B3A: data_out = 8'h95;
                    16'h5B3B: data_out = 8'h96;
                    16'h5B3C: data_out = 8'h97;
                    16'h5B3D: data_out = 8'h98;
                    16'h5B3E: data_out = 8'h99;
                    16'h5B3F: data_out = 8'h9A;
                    16'h5B40: data_out = 8'h9B;
                    16'h5B41: data_out = 8'h9C;
                    16'h5B42: data_out = 8'h9D;
                    16'h5B43: data_out = 8'h9E;
                    16'h5B44: data_out = 8'h9F;
                    16'h5B45: data_out = 8'hA0;
                    16'h5B46: data_out = 8'hA1;
                    16'h5B47: data_out = 8'hA2;
                    16'h5B48: data_out = 8'hA3;
                    16'h5B49: data_out = 8'hA4;
                    16'h5B4A: data_out = 8'hA5;
                    16'h5B4B: data_out = 8'hA6;
                    16'h5B4C: data_out = 8'hA7;
                    16'h5B4D: data_out = 8'hA8;
                    16'h5B4E: data_out = 8'hA9;
                    16'h5B4F: data_out = 8'hAA;
                    16'h5B50: data_out = 8'hAB;
                    16'h5B51: data_out = 8'hAC;
                    16'h5B52: data_out = 8'hAD;
                    16'h5B53: data_out = 8'hAE;
                    16'h5B54: data_out = 8'hAF;
                    16'h5B55: data_out = 8'hB0;
                    16'h5B56: data_out = 8'hB1;
                    16'h5B57: data_out = 8'hB2;
                    16'h5B58: data_out = 8'hB3;
                    16'h5B59: data_out = 8'hB4;
                    16'h5B5A: data_out = 8'hB5;
                    16'h5B5B: data_out = 8'hB6;
                    16'h5B5C: data_out = 8'hB7;
                    16'h5B5D: data_out = 8'hB8;
                    16'h5B5E: data_out = 8'hB9;
                    16'h5B5F: data_out = 8'hBA;
                    16'h5B60: data_out = 8'hBB;
                    16'h5B61: data_out = 8'hBC;
                    16'h5B62: data_out = 8'hBD;
                    16'h5B63: data_out = 8'hBE;
                    16'h5B64: data_out = 8'hBF;
                    16'h5B65: data_out = 8'hC0;
                    16'h5B66: data_out = 8'hC1;
                    16'h5B67: data_out = 8'hC2;
                    16'h5B68: data_out = 8'hC3;
                    16'h5B69: data_out = 8'hC4;
                    16'h5B6A: data_out = 8'hC5;
                    16'h5B6B: data_out = 8'hC6;
                    16'h5B6C: data_out = 8'hC7;
                    16'h5B6D: data_out = 8'hC8;
                    16'h5B6E: data_out = 8'hC9;
                    16'h5B6F: data_out = 8'hCA;
                    16'h5B70: data_out = 8'hCB;
                    16'h5B71: data_out = 8'hCC;
                    16'h5B72: data_out = 8'hCD;
                    16'h5B73: data_out = 8'hCE;
                    16'h5B74: data_out = 8'hCF;
                    16'h5B75: data_out = 8'hD0;
                    16'h5B76: data_out = 8'hD1;
                    16'h5B77: data_out = 8'hD2;
                    16'h5B78: data_out = 8'hD3;
                    16'h5B79: data_out = 8'hD4;
                    16'h5B7A: data_out = 8'hD5;
                    16'h5B7B: data_out = 8'hD6;
                    16'h5B7C: data_out = 8'hD7;
                    16'h5B7D: data_out = 8'hD8;
                    16'h5B7E: data_out = 8'hD9;
                    16'h5B7F: data_out = 8'hDA;
                    16'h5B80: data_out = 8'h5B;
                    16'h5B81: data_out = 8'h5A;
                    16'h5B82: data_out = 8'h59;
                    16'h5B83: data_out = 8'h58;
                    16'h5B84: data_out = 8'h57;
                    16'h5B85: data_out = 8'h56;
                    16'h5B86: data_out = 8'h55;
                    16'h5B87: data_out = 8'h54;
                    16'h5B88: data_out = 8'h53;
                    16'h5B89: data_out = 8'h52;
                    16'h5B8A: data_out = 8'h51;
                    16'h5B8B: data_out = 8'h50;
                    16'h5B8C: data_out = 8'h4F;
                    16'h5B8D: data_out = 8'h4E;
                    16'h5B8E: data_out = 8'h4D;
                    16'h5B8F: data_out = 8'h4C;
                    16'h5B90: data_out = 8'h4B;
                    16'h5B91: data_out = 8'h4A;
                    16'h5B92: data_out = 8'h49;
                    16'h5B93: data_out = 8'h48;
                    16'h5B94: data_out = 8'h47;
                    16'h5B95: data_out = 8'h46;
                    16'h5B96: data_out = 8'h45;
                    16'h5B97: data_out = 8'h44;
                    16'h5B98: data_out = 8'h43;
                    16'h5B99: data_out = 8'h42;
                    16'h5B9A: data_out = 8'h41;
                    16'h5B9B: data_out = 8'h40;
                    16'h5B9C: data_out = 8'h3F;
                    16'h5B9D: data_out = 8'h3E;
                    16'h5B9E: data_out = 8'h3D;
                    16'h5B9F: data_out = 8'h3C;
                    16'h5BA0: data_out = 8'h3B;
                    16'h5BA1: data_out = 8'h3A;
                    16'h5BA2: data_out = 8'h39;
                    16'h5BA3: data_out = 8'h38;
                    16'h5BA4: data_out = 8'h37;
                    16'h5BA5: data_out = 8'h36;
                    16'h5BA6: data_out = 8'h35;
                    16'h5BA7: data_out = 8'h34;
                    16'h5BA8: data_out = 8'h33;
                    16'h5BA9: data_out = 8'h32;
                    16'h5BAA: data_out = 8'h31;
                    16'h5BAB: data_out = 8'h30;
                    16'h5BAC: data_out = 8'h2F;
                    16'h5BAD: data_out = 8'h2E;
                    16'h5BAE: data_out = 8'h2D;
                    16'h5BAF: data_out = 8'h2C;
                    16'h5BB0: data_out = 8'h2B;
                    16'h5BB1: data_out = 8'h2A;
                    16'h5BB2: data_out = 8'h29;
                    16'h5BB3: data_out = 8'h28;
                    16'h5BB4: data_out = 8'h27;
                    16'h5BB5: data_out = 8'h26;
                    16'h5BB6: data_out = 8'h25;
                    16'h5BB7: data_out = 8'h24;
                    16'h5BB8: data_out = 8'h23;
                    16'h5BB9: data_out = 8'h22;
                    16'h5BBA: data_out = 8'h21;
                    16'h5BBB: data_out = 8'h20;
                    16'h5BBC: data_out = 8'h1F;
                    16'h5BBD: data_out = 8'h1E;
                    16'h5BBE: data_out = 8'h1D;
                    16'h5BBF: data_out = 8'h1C;
                    16'h5BC0: data_out = 8'h1B;
                    16'h5BC1: data_out = 8'h1A;
                    16'h5BC2: data_out = 8'h19;
                    16'h5BC3: data_out = 8'h18;
                    16'h5BC4: data_out = 8'h17;
                    16'h5BC5: data_out = 8'h16;
                    16'h5BC6: data_out = 8'h15;
                    16'h5BC7: data_out = 8'h14;
                    16'h5BC8: data_out = 8'h13;
                    16'h5BC9: data_out = 8'h12;
                    16'h5BCA: data_out = 8'h11;
                    16'h5BCB: data_out = 8'h10;
                    16'h5BCC: data_out = 8'hF;
                    16'h5BCD: data_out = 8'hE;
                    16'h5BCE: data_out = 8'hD;
                    16'h5BCF: data_out = 8'hC;
                    16'h5BD0: data_out = 8'hB;
                    16'h5BD1: data_out = 8'hA;
                    16'h5BD2: data_out = 8'h9;
                    16'h5BD3: data_out = 8'h8;
                    16'h5BD4: data_out = 8'h7;
                    16'h5BD5: data_out = 8'h6;
                    16'h5BD6: data_out = 8'h5;
                    16'h5BD7: data_out = 8'h4;
                    16'h5BD8: data_out = 8'h3;
                    16'h5BD9: data_out = 8'h2;
                    16'h5BDA: data_out = 8'h1;
                    16'h5BDB: data_out = 8'h0;
                    16'h5BDC: data_out = 8'h81;
                    16'h5BDD: data_out = 8'h82;
                    16'h5BDE: data_out = 8'h83;
                    16'h5BDF: data_out = 8'h84;
                    16'h5BE0: data_out = 8'h85;
                    16'h5BE1: data_out = 8'h86;
                    16'h5BE2: data_out = 8'h87;
                    16'h5BE3: data_out = 8'h88;
                    16'h5BE4: data_out = 8'h89;
                    16'h5BE5: data_out = 8'h8A;
                    16'h5BE6: data_out = 8'h8B;
                    16'h5BE7: data_out = 8'h8C;
                    16'h5BE8: data_out = 8'h8D;
                    16'h5BE9: data_out = 8'h8E;
                    16'h5BEA: data_out = 8'h8F;
                    16'h5BEB: data_out = 8'h90;
                    16'h5BEC: data_out = 8'h91;
                    16'h5BED: data_out = 8'h92;
                    16'h5BEE: data_out = 8'h93;
                    16'h5BEF: data_out = 8'h94;
                    16'h5BF0: data_out = 8'h95;
                    16'h5BF1: data_out = 8'h96;
                    16'h5BF2: data_out = 8'h97;
                    16'h5BF3: data_out = 8'h98;
                    16'h5BF4: data_out = 8'h99;
                    16'h5BF5: data_out = 8'h9A;
                    16'h5BF6: data_out = 8'h9B;
                    16'h5BF7: data_out = 8'h9C;
                    16'h5BF8: data_out = 8'h9D;
                    16'h5BF9: data_out = 8'h9E;
                    16'h5BFA: data_out = 8'h9F;
                    16'h5BFB: data_out = 8'hA0;
                    16'h5BFC: data_out = 8'hA1;
                    16'h5BFD: data_out = 8'hA2;
                    16'h5BFE: data_out = 8'hA3;
                    16'h5BFF: data_out = 8'hA4;
                    16'h5C00: data_out = 8'h5C;
                    16'h5C01: data_out = 8'h5D;
                    16'h5C02: data_out = 8'h5E;
                    16'h5C03: data_out = 8'h5F;
                    16'h5C04: data_out = 8'h60;
                    16'h5C05: data_out = 8'h61;
                    16'h5C06: data_out = 8'h62;
                    16'h5C07: data_out = 8'h63;
                    16'h5C08: data_out = 8'h64;
                    16'h5C09: data_out = 8'h65;
                    16'h5C0A: data_out = 8'h66;
                    16'h5C0B: data_out = 8'h67;
                    16'h5C0C: data_out = 8'h68;
                    16'h5C0D: data_out = 8'h69;
                    16'h5C0E: data_out = 8'h6A;
                    16'h5C0F: data_out = 8'h6B;
                    16'h5C10: data_out = 8'h6C;
                    16'h5C11: data_out = 8'h6D;
                    16'h5C12: data_out = 8'h6E;
                    16'h5C13: data_out = 8'h6F;
                    16'h5C14: data_out = 8'h70;
                    16'h5C15: data_out = 8'h71;
                    16'h5C16: data_out = 8'h72;
                    16'h5C17: data_out = 8'h73;
                    16'h5C18: data_out = 8'h74;
                    16'h5C19: data_out = 8'h75;
                    16'h5C1A: data_out = 8'h76;
                    16'h5C1B: data_out = 8'h77;
                    16'h5C1C: data_out = 8'h78;
                    16'h5C1D: data_out = 8'h79;
                    16'h5C1E: data_out = 8'h7A;
                    16'h5C1F: data_out = 8'h7B;
                    16'h5C20: data_out = 8'h7C;
                    16'h5C21: data_out = 8'h7D;
                    16'h5C22: data_out = 8'h7E;
                    16'h5C23: data_out = 8'h7F;
                    16'h5C24: data_out = 8'h80;
                    16'h5C25: data_out = 8'h81;
                    16'h5C26: data_out = 8'h82;
                    16'h5C27: data_out = 8'h83;
                    16'h5C28: data_out = 8'h84;
                    16'h5C29: data_out = 8'h85;
                    16'h5C2A: data_out = 8'h86;
                    16'h5C2B: data_out = 8'h87;
                    16'h5C2C: data_out = 8'h88;
                    16'h5C2D: data_out = 8'h89;
                    16'h5C2E: data_out = 8'h8A;
                    16'h5C2F: data_out = 8'h8B;
                    16'h5C30: data_out = 8'h8C;
                    16'h5C31: data_out = 8'h8D;
                    16'h5C32: data_out = 8'h8E;
                    16'h5C33: data_out = 8'h8F;
                    16'h5C34: data_out = 8'h90;
                    16'h5C35: data_out = 8'h91;
                    16'h5C36: data_out = 8'h92;
                    16'h5C37: data_out = 8'h93;
                    16'h5C38: data_out = 8'h94;
                    16'h5C39: data_out = 8'h95;
                    16'h5C3A: data_out = 8'h96;
                    16'h5C3B: data_out = 8'h97;
                    16'h5C3C: data_out = 8'h98;
                    16'h5C3D: data_out = 8'h99;
                    16'h5C3E: data_out = 8'h9A;
                    16'h5C3F: data_out = 8'h9B;
                    16'h5C40: data_out = 8'h9C;
                    16'h5C41: data_out = 8'h9D;
                    16'h5C42: data_out = 8'h9E;
                    16'h5C43: data_out = 8'h9F;
                    16'h5C44: data_out = 8'hA0;
                    16'h5C45: data_out = 8'hA1;
                    16'h5C46: data_out = 8'hA2;
                    16'h5C47: data_out = 8'hA3;
                    16'h5C48: data_out = 8'hA4;
                    16'h5C49: data_out = 8'hA5;
                    16'h5C4A: data_out = 8'hA6;
                    16'h5C4B: data_out = 8'hA7;
                    16'h5C4C: data_out = 8'hA8;
                    16'h5C4D: data_out = 8'hA9;
                    16'h5C4E: data_out = 8'hAA;
                    16'h5C4F: data_out = 8'hAB;
                    16'h5C50: data_out = 8'hAC;
                    16'h5C51: data_out = 8'hAD;
                    16'h5C52: data_out = 8'hAE;
                    16'h5C53: data_out = 8'hAF;
                    16'h5C54: data_out = 8'hB0;
                    16'h5C55: data_out = 8'hB1;
                    16'h5C56: data_out = 8'hB2;
                    16'h5C57: data_out = 8'hB3;
                    16'h5C58: data_out = 8'hB4;
                    16'h5C59: data_out = 8'hB5;
                    16'h5C5A: data_out = 8'hB6;
                    16'h5C5B: data_out = 8'hB7;
                    16'h5C5C: data_out = 8'hB8;
                    16'h5C5D: data_out = 8'hB9;
                    16'h5C5E: data_out = 8'hBA;
                    16'h5C5F: data_out = 8'hBB;
                    16'h5C60: data_out = 8'hBC;
                    16'h5C61: data_out = 8'hBD;
                    16'h5C62: data_out = 8'hBE;
                    16'h5C63: data_out = 8'hBF;
                    16'h5C64: data_out = 8'hC0;
                    16'h5C65: data_out = 8'hC1;
                    16'h5C66: data_out = 8'hC2;
                    16'h5C67: data_out = 8'hC3;
                    16'h5C68: data_out = 8'hC4;
                    16'h5C69: data_out = 8'hC5;
                    16'h5C6A: data_out = 8'hC6;
                    16'h5C6B: data_out = 8'hC7;
                    16'h5C6C: data_out = 8'hC8;
                    16'h5C6D: data_out = 8'hC9;
                    16'h5C6E: data_out = 8'hCA;
                    16'h5C6F: data_out = 8'hCB;
                    16'h5C70: data_out = 8'hCC;
                    16'h5C71: data_out = 8'hCD;
                    16'h5C72: data_out = 8'hCE;
                    16'h5C73: data_out = 8'hCF;
                    16'h5C74: data_out = 8'hD0;
                    16'h5C75: data_out = 8'hD1;
                    16'h5C76: data_out = 8'hD2;
                    16'h5C77: data_out = 8'hD3;
                    16'h5C78: data_out = 8'hD4;
                    16'h5C79: data_out = 8'hD5;
                    16'h5C7A: data_out = 8'hD6;
                    16'h5C7B: data_out = 8'hD7;
                    16'h5C7C: data_out = 8'hD8;
                    16'h5C7D: data_out = 8'hD9;
                    16'h5C7E: data_out = 8'hDA;
                    16'h5C7F: data_out = 8'hDB;
                    16'h5C80: data_out = 8'h5C;
                    16'h5C81: data_out = 8'h5B;
                    16'h5C82: data_out = 8'h5A;
                    16'h5C83: data_out = 8'h59;
                    16'h5C84: data_out = 8'h58;
                    16'h5C85: data_out = 8'h57;
                    16'h5C86: data_out = 8'h56;
                    16'h5C87: data_out = 8'h55;
                    16'h5C88: data_out = 8'h54;
                    16'h5C89: data_out = 8'h53;
                    16'h5C8A: data_out = 8'h52;
                    16'h5C8B: data_out = 8'h51;
                    16'h5C8C: data_out = 8'h50;
                    16'h5C8D: data_out = 8'h4F;
                    16'h5C8E: data_out = 8'h4E;
                    16'h5C8F: data_out = 8'h4D;
                    16'h5C90: data_out = 8'h4C;
                    16'h5C91: data_out = 8'h4B;
                    16'h5C92: data_out = 8'h4A;
                    16'h5C93: data_out = 8'h49;
                    16'h5C94: data_out = 8'h48;
                    16'h5C95: data_out = 8'h47;
                    16'h5C96: data_out = 8'h46;
                    16'h5C97: data_out = 8'h45;
                    16'h5C98: data_out = 8'h44;
                    16'h5C99: data_out = 8'h43;
                    16'h5C9A: data_out = 8'h42;
                    16'h5C9B: data_out = 8'h41;
                    16'h5C9C: data_out = 8'h40;
                    16'h5C9D: data_out = 8'h3F;
                    16'h5C9E: data_out = 8'h3E;
                    16'h5C9F: data_out = 8'h3D;
                    16'h5CA0: data_out = 8'h3C;
                    16'h5CA1: data_out = 8'h3B;
                    16'h5CA2: data_out = 8'h3A;
                    16'h5CA3: data_out = 8'h39;
                    16'h5CA4: data_out = 8'h38;
                    16'h5CA5: data_out = 8'h37;
                    16'h5CA6: data_out = 8'h36;
                    16'h5CA7: data_out = 8'h35;
                    16'h5CA8: data_out = 8'h34;
                    16'h5CA9: data_out = 8'h33;
                    16'h5CAA: data_out = 8'h32;
                    16'h5CAB: data_out = 8'h31;
                    16'h5CAC: data_out = 8'h30;
                    16'h5CAD: data_out = 8'h2F;
                    16'h5CAE: data_out = 8'h2E;
                    16'h5CAF: data_out = 8'h2D;
                    16'h5CB0: data_out = 8'h2C;
                    16'h5CB1: data_out = 8'h2B;
                    16'h5CB2: data_out = 8'h2A;
                    16'h5CB3: data_out = 8'h29;
                    16'h5CB4: data_out = 8'h28;
                    16'h5CB5: data_out = 8'h27;
                    16'h5CB6: data_out = 8'h26;
                    16'h5CB7: data_out = 8'h25;
                    16'h5CB8: data_out = 8'h24;
                    16'h5CB9: data_out = 8'h23;
                    16'h5CBA: data_out = 8'h22;
                    16'h5CBB: data_out = 8'h21;
                    16'h5CBC: data_out = 8'h20;
                    16'h5CBD: data_out = 8'h1F;
                    16'h5CBE: data_out = 8'h1E;
                    16'h5CBF: data_out = 8'h1D;
                    16'h5CC0: data_out = 8'h1C;
                    16'h5CC1: data_out = 8'h1B;
                    16'h5CC2: data_out = 8'h1A;
                    16'h5CC3: data_out = 8'h19;
                    16'h5CC4: data_out = 8'h18;
                    16'h5CC5: data_out = 8'h17;
                    16'h5CC6: data_out = 8'h16;
                    16'h5CC7: data_out = 8'h15;
                    16'h5CC8: data_out = 8'h14;
                    16'h5CC9: data_out = 8'h13;
                    16'h5CCA: data_out = 8'h12;
                    16'h5CCB: data_out = 8'h11;
                    16'h5CCC: data_out = 8'h10;
                    16'h5CCD: data_out = 8'hF;
                    16'h5CCE: data_out = 8'hE;
                    16'h5CCF: data_out = 8'hD;
                    16'h5CD0: data_out = 8'hC;
                    16'h5CD1: data_out = 8'hB;
                    16'h5CD2: data_out = 8'hA;
                    16'h5CD3: data_out = 8'h9;
                    16'h5CD4: data_out = 8'h8;
                    16'h5CD5: data_out = 8'h7;
                    16'h5CD6: data_out = 8'h6;
                    16'h5CD7: data_out = 8'h5;
                    16'h5CD8: data_out = 8'h4;
                    16'h5CD9: data_out = 8'h3;
                    16'h5CDA: data_out = 8'h2;
                    16'h5CDB: data_out = 8'h1;
                    16'h5CDC: data_out = 8'h0;
                    16'h5CDD: data_out = 8'h81;
                    16'h5CDE: data_out = 8'h82;
                    16'h5CDF: data_out = 8'h83;
                    16'h5CE0: data_out = 8'h84;
                    16'h5CE1: data_out = 8'h85;
                    16'h5CE2: data_out = 8'h86;
                    16'h5CE3: data_out = 8'h87;
                    16'h5CE4: data_out = 8'h88;
                    16'h5CE5: data_out = 8'h89;
                    16'h5CE6: data_out = 8'h8A;
                    16'h5CE7: data_out = 8'h8B;
                    16'h5CE8: data_out = 8'h8C;
                    16'h5CE9: data_out = 8'h8D;
                    16'h5CEA: data_out = 8'h8E;
                    16'h5CEB: data_out = 8'h8F;
                    16'h5CEC: data_out = 8'h90;
                    16'h5CED: data_out = 8'h91;
                    16'h5CEE: data_out = 8'h92;
                    16'h5CEF: data_out = 8'h93;
                    16'h5CF0: data_out = 8'h94;
                    16'h5CF1: data_out = 8'h95;
                    16'h5CF2: data_out = 8'h96;
                    16'h5CF3: data_out = 8'h97;
                    16'h5CF4: data_out = 8'h98;
                    16'h5CF5: data_out = 8'h99;
                    16'h5CF6: data_out = 8'h9A;
                    16'h5CF7: data_out = 8'h9B;
                    16'h5CF8: data_out = 8'h9C;
                    16'h5CF9: data_out = 8'h9D;
                    16'h5CFA: data_out = 8'h9E;
                    16'h5CFB: data_out = 8'h9F;
                    16'h5CFC: data_out = 8'hA0;
                    16'h5CFD: data_out = 8'hA1;
                    16'h5CFE: data_out = 8'hA2;
                    16'h5CFF: data_out = 8'hA3;
                    16'h5D00: data_out = 8'h5D;
                    16'h5D01: data_out = 8'h5E;
                    16'h5D02: data_out = 8'h5F;
                    16'h5D03: data_out = 8'h60;
                    16'h5D04: data_out = 8'h61;
                    16'h5D05: data_out = 8'h62;
                    16'h5D06: data_out = 8'h63;
                    16'h5D07: data_out = 8'h64;
                    16'h5D08: data_out = 8'h65;
                    16'h5D09: data_out = 8'h66;
                    16'h5D0A: data_out = 8'h67;
                    16'h5D0B: data_out = 8'h68;
                    16'h5D0C: data_out = 8'h69;
                    16'h5D0D: data_out = 8'h6A;
                    16'h5D0E: data_out = 8'h6B;
                    16'h5D0F: data_out = 8'h6C;
                    16'h5D10: data_out = 8'h6D;
                    16'h5D11: data_out = 8'h6E;
                    16'h5D12: data_out = 8'h6F;
                    16'h5D13: data_out = 8'h70;
                    16'h5D14: data_out = 8'h71;
                    16'h5D15: data_out = 8'h72;
                    16'h5D16: data_out = 8'h73;
                    16'h5D17: data_out = 8'h74;
                    16'h5D18: data_out = 8'h75;
                    16'h5D19: data_out = 8'h76;
                    16'h5D1A: data_out = 8'h77;
                    16'h5D1B: data_out = 8'h78;
                    16'h5D1C: data_out = 8'h79;
                    16'h5D1D: data_out = 8'h7A;
                    16'h5D1E: data_out = 8'h7B;
                    16'h5D1F: data_out = 8'h7C;
                    16'h5D20: data_out = 8'h7D;
                    16'h5D21: data_out = 8'h7E;
                    16'h5D22: data_out = 8'h7F;
                    16'h5D23: data_out = 8'h80;
                    16'h5D24: data_out = 8'h81;
                    16'h5D25: data_out = 8'h82;
                    16'h5D26: data_out = 8'h83;
                    16'h5D27: data_out = 8'h84;
                    16'h5D28: data_out = 8'h85;
                    16'h5D29: data_out = 8'h86;
                    16'h5D2A: data_out = 8'h87;
                    16'h5D2B: data_out = 8'h88;
                    16'h5D2C: data_out = 8'h89;
                    16'h5D2D: data_out = 8'h8A;
                    16'h5D2E: data_out = 8'h8B;
                    16'h5D2F: data_out = 8'h8C;
                    16'h5D30: data_out = 8'h8D;
                    16'h5D31: data_out = 8'h8E;
                    16'h5D32: data_out = 8'h8F;
                    16'h5D33: data_out = 8'h90;
                    16'h5D34: data_out = 8'h91;
                    16'h5D35: data_out = 8'h92;
                    16'h5D36: data_out = 8'h93;
                    16'h5D37: data_out = 8'h94;
                    16'h5D38: data_out = 8'h95;
                    16'h5D39: data_out = 8'h96;
                    16'h5D3A: data_out = 8'h97;
                    16'h5D3B: data_out = 8'h98;
                    16'h5D3C: data_out = 8'h99;
                    16'h5D3D: data_out = 8'h9A;
                    16'h5D3E: data_out = 8'h9B;
                    16'h5D3F: data_out = 8'h9C;
                    16'h5D40: data_out = 8'h9D;
                    16'h5D41: data_out = 8'h9E;
                    16'h5D42: data_out = 8'h9F;
                    16'h5D43: data_out = 8'hA0;
                    16'h5D44: data_out = 8'hA1;
                    16'h5D45: data_out = 8'hA2;
                    16'h5D46: data_out = 8'hA3;
                    16'h5D47: data_out = 8'hA4;
                    16'h5D48: data_out = 8'hA5;
                    16'h5D49: data_out = 8'hA6;
                    16'h5D4A: data_out = 8'hA7;
                    16'h5D4B: data_out = 8'hA8;
                    16'h5D4C: data_out = 8'hA9;
                    16'h5D4D: data_out = 8'hAA;
                    16'h5D4E: data_out = 8'hAB;
                    16'h5D4F: data_out = 8'hAC;
                    16'h5D50: data_out = 8'hAD;
                    16'h5D51: data_out = 8'hAE;
                    16'h5D52: data_out = 8'hAF;
                    16'h5D53: data_out = 8'hB0;
                    16'h5D54: data_out = 8'hB1;
                    16'h5D55: data_out = 8'hB2;
                    16'h5D56: data_out = 8'hB3;
                    16'h5D57: data_out = 8'hB4;
                    16'h5D58: data_out = 8'hB5;
                    16'h5D59: data_out = 8'hB6;
                    16'h5D5A: data_out = 8'hB7;
                    16'h5D5B: data_out = 8'hB8;
                    16'h5D5C: data_out = 8'hB9;
                    16'h5D5D: data_out = 8'hBA;
                    16'h5D5E: data_out = 8'hBB;
                    16'h5D5F: data_out = 8'hBC;
                    16'h5D60: data_out = 8'hBD;
                    16'h5D61: data_out = 8'hBE;
                    16'h5D62: data_out = 8'hBF;
                    16'h5D63: data_out = 8'hC0;
                    16'h5D64: data_out = 8'hC1;
                    16'h5D65: data_out = 8'hC2;
                    16'h5D66: data_out = 8'hC3;
                    16'h5D67: data_out = 8'hC4;
                    16'h5D68: data_out = 8'hC5;
                    16'h5D69: data_out = 8'hC6;
                    16'h5D6A: data_out = 8'hC7;
                    16'h5D6B: data_out = 8'hC8;
                    16'h5D6C: data_out = 8'hC9;
                    16'h5D6D: data_out = 8'hCA;
                    16'h5D6E: data_out = 8'hCB;
                    16'h5D6F: data_out = 8'hCC;
                    16'h5D70: data_out = 8'hCD;
                    16'h5D71: data_out = 8'hCE;
                    16'h5D72: data_out = 8'hCF;
                    16'h5D73: data_out = 8'hD0;
                    16'h5D74: data_out = 8'hD1;
                    16'h5D75: data_out = 8'hD2;
                    16'h5D76: data_out = 8'hD3;
                    16'h5D77: data_out = 8'hD4;
                    16'h5D78: data_out = 8'hD5;
                    16'h5D79: data_out = 8'hD6;
                    16'h5D7A: data_out = 8'hD7;
                    16'h5D7B: data_out = 8'hD8;
                    16'h5D7C: data_out = 8'hD9;
                    16'h5D7D: data_out = 8'hDA;
                    16'h5D7E: data_out = 8'hDB;
                    16'h5D7F: data_out = 8'hDC;
                    16'h5D80: data_out = 8'h5D;
                    16'h5D81: data_out = 8'h5C;
                    16'h5D82: data_out = 8'h5B;
                    16'h5D83: data_out = 8'h5A;
                    16'h5D84: data_out = 8'h59;
                    16'h5D85: data_out = 8'h58;
                    16'h5D86: data_out = 8'h57;
                    16'h5D87: data_out = 8'h56;
                    16'h5D88: data_out = 8'h55;
                    16'h5D89: data_out = 8'h54;
                    16'h5D8A: data_out = 8'h53;
                    16'h5D8B: data_out = 8'h52;
                    16'h5D8C: data_out = 8'h51;
                    16'h5D8D: data_out = 8'h50;
                    16'h5D8E: data_out = 8'h4F;
                    16'h5D8F: data_out = 8'h4E;
                    16'h5D90: data_out = 8'h4D;
                    16'h5D91: data_out = 8'h4C;
                    16'h5D92: data_out = 8'h4B;
                    16'h5D93: data_out = 8'h4A;
                    16'h5D94: data_out = 8'h49;
                    16'h5D95: data_out = 8'h48;
                    16'h5D96: data_out = 8'h47;
                    16'h5D97: data_out = 8'h46;
                    16'h5D98: data_out = 8'h45;
                    16'h5D99: data_out = 8'h44;
                    16'h5D9A: data_out = 8'h43;
                    16'h5D9B: data_out = 8'h42;
                    16'h5D9C: data_out = 8'h41;
                    16'h5D9D: data_out = 8'h40;
                    16'h5D9E: data_out = 8'h3F;
                    16'h5D9F: data_out = 8'h3E;
                    16'h5DA0: data_out = 8'h3D;
                    16'h5DA1: data_out = 8'h3C;
                    16'h5DA2: data_out = 8'h3B;
                    16'h5DA3: data_out = 8'h3A;
                    16'h5DA4: data_out = 8'h39;
                    16'h5DA5: data_out = 8'h38;
                    16'h5DA6: data_out = 8'h37;
                    16'h5DA7: data_out = 8'h36;
                    16'h5DA8: data_out = 8'h35;
                    16'h5DA9: data_out = 8'h34;
                    16'h5DAA: data_out = 8'h33;
                    16'h5DAB: data_out = 8'h32;
                    16'h5DAC: data_out = 8'h31;
                    16'h5DAD: data_out = 8'h30;
                    16'h5DAE: data_out = 8'h2F;
                    16'h5DAF: data_out = 8'h2E;
                    16'h5DB0: data_out = 8'h2D;
                    16'h5DB1: data_out = 8'h2C;
                    16'h5DB2: data_out = 8'h2B;
                    16'h5DB3: data_out = 8'h2A;
                    16'h5DB4: data_out = 8'h29;
                    16'h5DB5: data_out = 8'h28;
                    16'h5DB6: data_out = 8'h27;
                    16'h5DB7: data_out = 8'h26;
                    16'h5DB8: data_out = 8'h25;
                    16'h5DB9: data_out = 8'h24;
                    16'h5DBA: data_out = 8'h23;
                    16'h5DBB: data_out = 8'h22;
                    16'h5DBC: data_out = 8'h21;
                    16'h5DBD: data_out = 8'h20;
                    16'h5DBE: data_out = 8'h1F;
                    16'h5DBF: data_out = 8'h1E;
                    16'h5DC0: data_out = 8'h1D;
                    16'h5DC1: data_out = 8'h1C;
                    16'h5DC2: data_out = 8'h1B;
                    16'h5DC3: data_out = 8'h1A;
                    16'h5DC4: data_out = 8'h19;
                    16'h5DC5: data_out = 8'h18;
                    16'h5DC6: data_out = 8'h17;
                    16'h5DC7: data_out = 8'h16;
                    16'h5DC8: data_out = 8'h15;
                    16'h5DC9: data_out = 8'h14;
                    16'h5DCA: data_out = 8'h13;
                    16'h5DCB: data_out = 8'h12;
                    16'h5DCC: data_out = 8'h11;
                    16'h5DCD: data_out = 8'h10;
                    16'h5DCE: data_out = 8'hF;
                    16'h5DCF: data_out = 8'hE;
                    16'h5DD0: data_out = 8'hD;
                    16'h5DD1: data_out = 8'hC;
                    16'h5DD2: data_out = 8'hB;
                    16'h5DD3: data_out = 8'hA;
                    16'h5DD4: data_out = 8'h9;
                    16'h5DD5: data_out = 8'h8;
                    16'h5DD6: data_out = 8'h7;
                    16'h5DD7: data_out = 8'h6;
                    16'h5DD8: data_out = 8'h5;
                    16'h5DD9: data_out = 8'h4;
                    16'h5DDA: data_out = 8'h3;
                    16'h5DDB: data_out = 8'h2;
                    16'h5DDC: data_out = 8'h1;
                    16'h5DDD: data_out = 8'h0;
                    16'h5DDE: data_out = 8'h81;
                    16'h5DDF: data_out = 8'h82;
                    16'h5DE0: data_out = 8'h83;
                    16'h5DE1: data_out = 8'h84;
                    16'h5DE2: data_out = 8'h85;
                    16'h5DE3: data_out = 8'h86;
                    16'h5DE4: data_out = 8'h87;
                    16'h5DE5: data_out = 8'h88;
                    16'h5DE6: data_out = 8'h89;
                    16'h5DE7: data_out = 8'h8A;
                    16'h5DE8: data_out = 8'h8B;
                    16'h5DE9: data_out = 8'h8C;
                    16'h5DEA: data_out = 8'h8D;
                    16'h5DEB: data_out = 8'h8E;
                    16'h5DEC: data_out = 8'h8F;
                    16'h5DED: data_out = 8'h90;
                    16'h5DEE: data_out = 8'h91;
                    16'h5DEF: data_out = 8'h92;
                    16'h5DF0: data_out = 8'h93;
                    16'h5DF1: data_out = 8'h94;
                    16'h5DF2: data_out = 8'h95;
                    16'h5DF3: data_out = 8'h96;
                    16'h5DF4: data_out = 8'h97;
                    16'h5DF5: data_out = 8'h98;
                    16'h5DF6: data_out = 8'h99;
                    16'h5DF7: data_out = 8'h9A;
                    16'h5DF8: data_out = 8'h9B;
                    16'h5DF9: data_out = 8'h9C;
                    16'h5DFA: data_out = 8'h9D;
                    16'h5DFB: data_out = 8'h9E;
                    16'h5DFC: data_out = 8'h9F;
                    16'h5DFD: data_out = 8'hA0;
                    16'h5DFE: data_out = 8'hA1;
                    16'h5DFF: data_out = 8'hA2;
                    16'h5E00: data_out = 8'h5E;
                    16'h5E01: data_out = 8'h5F;
                    16'h5E02: data_out = 8'h60;
                    16'h5E03: data_out = 8'h61;
                    16'h5E04: data_out = 8'h62;
                    16'h5E05: data_out = 8'h63;
                    16'h5E06: data_out = 8'h64;
                    16'h5E07: data_out = 8'h65;
                    16'h5E08: data_out = 8'h66;
                    16'h5E09: data_out = 8'h67;
                    16'h5E0A: data_out = 8'h68;
                    16'h5E0B: data_out = 8'h69;
                    16'h5E0C: data_out = 8'h6A;
                    16'h5E0D: data_out = 8'h6B;
                    16'h5E0E: data_out = 8'h6C;
                    16'h5E0F: data_out = 8'h6D;
                    16'h5E10: data_out = 8'h6E;
                    16'h5E11: data_out = 8'h6F;
                    16'h5E12: data_out = 8'h70;
                    16'h5E13: data_out = 8'h71;
                    16'h5E14: data_out = 8'h72;
                    16'h5E15: data_out = 8'h73;
                    16'h5E16: data_out = 8'h74;
                    16'h5E17: data_out = 8'h75;
                    16'h5E18: data_out = 8'h76;
                    16'h5E19: data_out = 8'h77;
                    16'h5E1A: data_out = 8'h78;
                    16'h5E1B: data_out = 8'h79;
                    16'h5E1C: data_out = 8'h7A;
                    16'h5E1D: data_out = 8'h7B;
                    16'h5E1E: data_out = 8'h7C;
                    16'h5E1F: data_out = 8'h7D;
                    16'h5E20: data_out = 8'h7E;
                    16'h5E21: data_out = 8'h7F;
                    16'h5E22: data_out = 8'h80;
                    16'h5E23: data_out = 8'h81;
                    16'h5E24: data_out = 8'h82;
                    16'h5E25: data_out = 8'h83;
                    16'h5E26: data_out = 8'h84;
                    16'h5E27: data_out = 8'h85;
                    16'h5E28: data_out = 8'h86;
                    16'h5E29: data_out = 8'h87;
                    16'h5E2A: data_out = 8'h88;
                    16'h5E2B: data_out = 8'h89;
                    16'h5E2C: data_out = 8'h8A;
                    16'h5E2D: data_out = 8'h8B;
                    16'h5E2E: data_out = 8'h8C;
                    16'h5E2F: data_out = 8'h8D;
                    16'h5E30: data_out = 8'h8E;
                    16'h5E31: data_out = 8'h8F;
                    16'h5E32: data_out = 8'h90;
                    16'h5E33: data_out = 8'h91;
                    16'h5E34: data_out = 8'h92;
                    16'h5E35: data_out = 8'h93;
                    16'h5E36: data_out = 8'h94;
                    16'h5E37: data_out = 8'h95;
                    16'h5E38: data_out = 8'h96;
                    16'h5E39: data_out = 8'h97;
                    16'h5E3A: data_out = 8'h98;
                    16'h5E3B: data_out = 8'h99;
                    16'h5E3C: data_out = 8'h9A;
                    16'h5E3D: data_out = 8'h9B;
                    16'h5E3E: data_out = 8'h9C;
                    16'h5E3F: data_out = 8'h9D;
                    16'h5E40: data_out = 8'h9E;
                    16'h5E41: data_out = 8'h9F;
                    16'h5E42: data_out = 8'hA0;
                    16'h5E43: data_out = 8'hA1;
                    16'h5E44: data_out = 8'hA2;
                    16'h5E45: data_out = 8'hA3;
                    16'h5E46: data_out = 8'hA4;
                    16'h5E47: data_out = 8'hA5;
                    16'h5E48: data_out = 8'hA6;
                    16'h5E49: data_out = 8'hA7;
                    16'h5E4A: data_out = 8'hA8;
                    16'h5E4B: data_out = 8'hA9;
                    16'h5E4C: data_out = 8'hAA;
                    16'h5E4D: data_out = 8'hAB;
                    16'h5E4E: data_out = 8'hAC;
                    16'h5E4F: data_out = 8'hAD;
                    16'h5E50: data_out = 8'hAE;
                    16'h5E51: data_out = 8'hAF;
                    16'h5E52: data_out = 8'hB0;
                    16'h5E53: data_out = 8'hB1;
                    16'h5E54: data_out = 8'hB2;
                    16'h5E55: data_out = 8'hB3;
                    16'h5E56: data_out = 8'hB4;
                    16'h5E57: data_out = 8'hB5;
                    16'h5E58: data_out = 8'hB6;
                    16'h5E59: data_out = 8'hB7;
                    16'h5E5A: data_out = 8'hB8;
                    16'h5E5B: data_out = 8'hB9;
                    16'h5E5C: data_out = 8'hBA;
                    16'h5E5D: data_out = 8'hBB;
                    16'h5E5E: data_out = 8'hBC;
                    16'h5E5F: data_out = 8'hBD;
                    16'h5E60: data_out = 8'hBE;
                    16'h5E61: data_out = 8'hBF;
                    16'h5E62: data_out = 8'hC0;
                    16'h5E63: data_out = 8'hC1;
                    16'h5E64: data_out = 8'hC2;
                    16'h5E65: data_out = 8'hC3;
                    16'h5E66: data_out = 8'hC4;
                    16'h5E67: data_out = 8'hC5;
                    16'h5E68: data_out = 8'hC6;
                    16'h5E69: data_out = 8'hC7;
                    16'h5E6A: data_out = 8'hC8;
                    16'h5E6B: data_out = 8'hC9;
                    16'h5E6C: data_out = 8'hCA;
                    16'h5E6D: data_out = 8'hCB;
                    16'h5E6E: data_out = 8'hCC;
                    16'h5E6F: data_out = 8'hCD;
                    16'h5E70: data_out = 8'hCE;
                    16'h5E71: data_out = 8'hCF;
                    16'h5E72: data_out = 8'hD0;
                    16'h5E73: data_out = 8'hD1;
                    16'h5E74: data_out = 8'hD2;
                    16'h5E75: data_out = 8'hD3;
                    16'h5E76: data_out = 8'hD4;
                    16'h5E77: data_out = 8'hD5;
                    16'h5E78: data_out = 8'hD6;
                    16'h5E79: data_out = 8'hD7;
                    16'h5E7A: data_out = 8'hD8;
                    16'h5E7B: data_out = 8'hD9;
                    16'h5E7C: data_out = 8'hDA;
                    16'h5E7D: data_out = 8'hDB;
                    16'h5E7E: data_out = 8'hDC;
                    16'h5E7F: data_out = 8'hDD;
                    16'h5E80: data_out = 8'h5E;
                    16'h5E81: data_out = 8'h5D;
                    16'h5E82: data_out = 8'h5C;
                    16'h5E83: data_out = 8'h5B;
                    16'h5E84: data_out = 8'h5A;
                    16'h5E85: data_out = 8'h59;
                    16'h5E86: data_out = 8'h58;
                    16'h5E87: data_out = 8'h57;
                    16'h5E88: data_out = 8'h56;
                    16'h5E89: data_out = 8'h55;
                    16'h5E8A: data_out = 8'h54;
                    16'h5E8B: data_out = 8'h53;
                    16'h5E8C: data_out = 8'h52;
                    16'h5E8D: data_out = 8'h51;
                    16'h5E8E: data_out = 8'h50;
                    16'h5E8F: data_out = 8'h4F;
                    16'h5E90: data_out = 8'h4E;
                    16'h5E91: data_out = 8'h4D;
                    16'h5E92: data_out = 8'h4C;
                    16'h5E93: data_out = 8'h4B;
                    16'h5E94: data_out = 8'h4A;
                    16'h5E95: data_out = 8'h49;
                    16'h5E96: data_out = 8'h48;
                    16'h5E97: data_out = 8'h47;
                    16'h5E98: data_out = 8'h46;
                    16'h5E99: data_out = 8'h45;
                    16'h5E9A: data_out = 8'h44;
                    16'h5E9B: data_out = 8'h43;
                    16'h5E9C: data_out = 8'h42;
                    16'h5E9D: data_out = 8'h41;
                    16'h5E9E: data_out = 8'h40;
                    16'h5E9F: data_out = 8'h3F;
                    16'h5EA0: data_out = 8'h3E;
                    16'h5EA1: data_out = 8'h3D;
                    16'h5EA2: data_out = 8'h3C;
                    16'h5EA3: data_out = 8'h3B;
                    16'h5EA4: data_out = 8'h3A;
                    16'h5EA5: data_out = 8'h39;
                    16'h5EA6: data_out = 8'h38;
                    16'h5EA7: data_out = 8'h37;
                    16'h5EA8: data_out = 8'h36;
                    16'h5EA9: data_out = 8'h35;
                    16'h5EAA: data_out = 8'h34;
                    16'h5EAB: data_out = 8'h33;
                    16'h5EAC: data_out = 8'h32;
                    16'h5EAD: data_out = 8'h31;
                    16'h5EAE: data_out = 8'h30;
                    16'h5EAF: data_out = 8'h2F;
                    16'h5EB0: data_out = 8'h2E;
                    16'h5EB1: data_out = 8'h2D;
                    16'h5EB2: data_out = 8'h2C;
                    16'h5EB3: data_out = 8'h2B;
                    16'h5EB4: data_out = 8'h2A;
                    16'h5EB5: data_out = 8'h29;
                    16'h5EB6: data_out = 8'h28;
                    16'h5EB7: data_out = 8'h27;
                    16'h5EB8: data_out = 8'h26;
                    16'h5EB9: data_out = 8'h25;
                    16'h5EBA: data_out = 8'h24;
                    16'h5EBB: data_out = 8'h23;
                    16'h5EBC: data_out = 8'h22;
                    16'h5EBD: data_out = 8'h21;
                    16'h5EBE: data_out = 8'h20;
                    16'h5EBF: data_out = 8'h1F;
                    16'h5EC0: data_out = 8'h1E;
                    16'h5EC1: data_out = 8'h1D;
                    16'h5EC2: data_out = 8'h1C;
                    16'h5EC3: data_out = 8'h1B;
                    16'h5EC4: data_out = 8'h1A;
                    16'h5EC5: data_out = 8'h19;
                    16'h5EC6: data_out = 8'h18;
                    16'h5EC7: data_out = 8'h17;
                    16'h5EC8: data_out = 8'h16;
                    16'h5EC9: data_out = 8'h15;
                    16'h5ECA: data_out = 8'h14;
                    16'h5ECB: data_out = 8'h13;
                    16'h5ECC: data_out = 8'h12;
                    16'h5ECD: data_out = 8'h11;
                    16'h5ECE: data_out = 8'h10;
                    16'h5ECF: data_out = 8'hF;
                    16'h5ED0: data_out = 8'hE;
                    16'h5ED1: data_out = 8'hD;
                    16'h5ED2: data_out = 8'hC;
                    16'h5ED3: data_out = 8'hB;
                    16'h5ED4: data_out = 8'hA;
                    16'h5ED5: data_out = 8'h9;
                    16'h5ED6: data_out = 8'h8;
                    16'h5ED7: data_out = 8'h7;
                    16'h5ED8: data_out = 8'h6;
                    16'h5ED9: data_out = 8'h5;
                    16'h5EDA: data_out = 8'h4;
                    16'h5EDB: data_out = 8'h3;
                    16'h5EDC: data_out = 8'h2;
                    16'h5EDD: data_out = 8'h1;
                    16'h5EDE: data_out = 8'h0;
                    16'h5EDF: data_out = 8'h81;
                    16'h5EE0: data_out = 8'h82;
                    16'h5EE1: data_out = 8'h83;
                    16'h5EE2: data_out = 8'h84;
                    16'h5EE3: data_out = 8'h85;
                    16'h5EE4: data_out = 8'h86;
                    16'h5EE5: data_out = 8'h87;
                    16'h5EE6: data_out = 8'h88;
                    16'h5EE7: data_out = 8'h89;
                    16'h5EE8: data_out = 8'h8A;
                    16'h5EE9: data_out = 8'h8B;
                    16'h5EEA: data_out = 8'h8C;
                    16'h5EEB: data_out = 8'h8D;
                    16'h5EEC: data_out = 8'h8E;
                    16'h5EED: data_out = 8'h8F;
                    16'h5EEE: data_out = 8'h90;
                    16'h5EEF: data_out = 8'h91;
                    16'h5EF0: data_out = 8'h92;
                    16'h5EF1: data_out = 8'h93;
                    16'h5EF2: data_out = 8'h94;
                    16'h5EF3: data_out = 8'h95;
                    16'h5EF4: data_out = 8'h96;
                    16'h5EF5: data_out = 8'h97;
                    16'h5EF6: data_out = 8'h98;
                    16'h5EF7: data_out = 8'h99;
                    16'h5EF8: data_out = 8'h9A;
                    16'h5EF9: data_out = 8'h9B;
                    16'h5EFA: data_out = 8'h9C;
                    16'h5EFB: data_out = 8'h9D;
                    16'h5EFC: data_out = 8'h9E;
                    16'h5EFD: data_out = 8'h9F;
                    16'h5EFE: data_out = 8'hA0;
                    16'h5EFF: data_out = 8'hA1;
                    16'h5F00: data_out = 8'h5F;
                    16'h5F01: data_out = 8'h60;
                    16'h5F02: data_out = 8'h61;
                    16'h5F03: data_out = 8'h62;
                    16'h5F04: data_out = 8'h63;
                    16'h5F05: data_out = 8'h64;
                    16'h5F06: data_out = 8'h65;
                    16'h5F07: data_out = 8'h66;
                    16'h5F08: data_out = 8'h67;
                    16'h5F09: data_out = 8'h68;
                    16'h5F0A: data_out = 8'h69;
                    16'h5F0B: data_out = 8'h6A;
                    16'h5F0C: data_out = 8'h6B;
                    16'h5F0D: data_out = 8'h6C;
                    16'h5F0E: data_out = 8'h6D;
                    16'h5F0F: data_out = 8'h6E;
                    16'h5F10: data_out = 8'h6F;
                    16'h5F11: data_out = 8'h70;
                    16'h5F12: data_out = 8'h71;
                    16'h5F13: data_out = 8'h72;
                    16'h5F14: data_out = 8'h73;
                    16'h5F15: data_out = 8'h74;
                    16'h5F16: data_out = 8'h75;
                    16'h5F17: data_out = 8'h76;
                    16'h5F18: data_out = 8'h77;
                    16'h5F19: data_out = 8'h78;
                    16'h5F1A: data_out = 8'h79;
                    16'h5F1B: data_out = 8'h7A;
                    16'h5F1C: data_out = 8'h7B;
                    16'h5F1D: data_out = 8'h7C;
                    16'h5F1E: data_out = 8'h7D;
                    16'h5F1F: data_out = 8'h7E;
                    16'h5F20: data_out = 8'h7F;
                    16'h5F21: data_out = 8'h80;
                    16'h5F22: data_out = 8'h81;
                    16'h5F23: data_out = 8'h82;
                    16'h5F24: data_out = 8'h83;
                    16'h5F25: data_out = 8'h84;
                    16'h5F26: data_out = 8'h85;
                    16'h5F27: data_out = 8'h86;
                    16'h5F28: data_out = 8'h87;
                    16'h5F29: data_out = 8'h88;
                    16'h5F2A: data_out = 8'h89;
                    16'h5F2B: data_out = 8'h8A;
                    16'h5F2C: data_out = 8'h8B;
                    16'h5F2D: data_out = 8'h8C;
                    16'h5F2E: data_out = 8'h8D;
                    16'h5F2F: data_out = 8'h8E;
                    16'h5F30: data_out = 8'h8F;
                    16'h5F31: data_out = 8'h90;
                    16'h5F32: data_out = 8'h91;
                    16'h5F33: data_out = 8'h92;
                    16'h5F34: data_out = 8'h93;
                    16'h5F35: data_out = 8'h94;
                    16'h5F36: data_out = 8'h95;
                    16'h5F37: data_out = 8'h96;
                    16'h5F38: data_out = 8'h97;
                    16'h5F39: data_out = 8'h98;
                    16'h5F3A: data_out = 8'h99;
                    16'h5F3B: data_out = 8'h9A;
                    16'h5F3C: data_out = 8'h9B;
                    16'h5F3D: data_out = 8'h9C;
                    16'h5F3E: data_out = 8'h9D;
                    16'h5F3F: data_out = 8'h9E;
                    16'h5F40: data_out = 8'h9F;
                    16'h5F41: data_out = 8'hA0;
                    16'h5F42: data_out = 8'hA1;
                    16'h5F43: data_out = 8'hA2;
                    16'h5F44: data_out = 8'hA3;
                    16'h5F45: data_out = 8'hA4;
                    16'h5F46: data_out = 8'hA5;
                    16'h5F47: data_out = 8'hA6;
                    16'h5F48: data_out = 8'hA7;
                    16'h5F49: data_out = 8'hA8;
                    16'h5F4A: data_out = 8'hA9;
                    16'h5F4B: data_out = 8'hAA;
                    16'h5F4C: data_out = 8'hAB;
                    16'h5F4D: data_out = 8'hAC;
                    16'h5F4E: data_out = 8'hAD;
                    16'h5F4F: data_out = 8'hAE;
                    16'h5F50: data_out = 8'hAF;
                    16'h5F51: data_out = 8'hB0;
                    16'h5F52: data_out = 8'hB1;
                    16'h5F53: data_out = 8'hB2;
                    16'h5F54: data_out = 8'hB3;
                    16'h5F55: data_out = 8'hB4;
                    16'h5F56: data_out = 8'hB5;
                    16'h5F57: data_out = 8'hB6;
                    16'h5F58: data_out = 8'hB7;
                    16'h5F59: data_out = 8'hB8;
                    16'h5F5A: data_out = 8'hB9;
                    16'h5F5B: data_out = 8'hBA;
                    16'h5F5C: data_out = 8'hBB;
                    16'h5F5D: data_out = 8'hBC;
                    16'h5F5E: data_out = 8'hBD;
                    16'h5F5F: data_out = 8'hBE;
                    16'h5F60: data_out = 8'hBF;
                    16'h5F61: data_out = 8'hC0;
                    16'h5F62: data_out = 8'hC1;
                    16'h5F63: data_out = 8'hC2;
                    16'h5F64: data_out = 8'hC3;
                    16'h5F65: data_out = 8'hC4;
                    16'h5F66: data_out = 8'hC5;
                    16'h5F67: data_out = 8'hC6;
                    16'h5F68: data_out = 8'hC7;
                    16'h5F69: data_out = 8'hC8;
                    16'h5F6A: data_out = 8'hC9;
                    16'h5F6B: data_out = 8'hCA;
                    16'h5F6C: data_out = 8'hCB;
                    16'h5F6D: data_out = 8'hCC;
                    16'h5F6E: data_out = 8'hCD;
                    16'h5F6F: data_out = 8'hCE;
                    16'h5F70: data_out = 8'hCF;
                    16'h5F71: data_out = 8'hD0;
                    16'h5F72: data_out = 8'hD1;
                    16'h5F73: data_out = 8'hD2;
                    16'h5F74: data_out = 8'hD3;
                    16'h5F75: data_out = 8'hD4;
                    16'h5F76: data_out = 8'hD5;
                    16'h5F77: data_out = 8'hD6;
                    16'h5F78: data_out = 8'hD7;
                    16'h5F79: data_out = 8'hD8;
                    16'h5F7A: data_out = 8'hD9;
                    16'h5F7B: data_out = 8'hDA;
                    16'h5F7C: data_out = 8'hDB;
                    16'h5F7D: data_out = 8'hDC;
                    16'h5F7E: data_out = 8'hDD;
                    16'h5F7F: data_out = 8'hDE;
                    16'h5F80: data_out = 8'h5F;
                    16'h5F81: data_out = 8'h5E;
                    16'h5F82: data_out = 8'h5D;
                    16'h5F83: data_out = 8'h5C;
                    16'h5F84: data_out = 8'h5B;
                    16'h5F85: data_out = 8'h5A;
                    16'h5F86: data_out = 8'h59;
                    16'h5F87: data_out = 8'h58;
                    16'h5F88: data_out = 8'h57;
                    16'h5F89: data_out = 8'h56;
                    16'h5F8A: data_out = 8'h55;
                    16'h5F8B: data_out = 8'h54;
                    16'h5F8C: data_out = 8'h53;
                    16'h5F8D: data_out = 8'h52;
                    16'h5F8E: data_out = 8'h51;
                    16'h5F8F: data_out = 8'h50;
                    16'h5F90: data_out = 8'h4F;
                    16'h5F91: data_out = 8'h4E;
                    16'h5F92: data_out = 8'h4D;
                    16'h5F93: data_out = 8'h4C;
                    16'h5F94: data_out = 8'h4B;
                    16'h5F95: data_out = 8'h4A;
                    16'h5F96: data_out = 8'h49;
                    16'h5F97: data_out = 8'h48;
                    16'h5F98: data_out = 8'h47;
                    16'h5F99: data_out = 8'h46;
                    16'h5F9A: data_out = 8'h45;
                    16'h5F9B: data_out = 8'h44;
                    16'h5F9C: data_out = 8'h43;
                    16'h5F9D: data_out = 8'h42;
                    16'h5F9E: data_out = 8'h41;
                    16'h5F9F: data_out = 8'h40;
                    16'h5FA0: data_out = 8'h3F;
                    16'h5FA1: data_out = 8'h3E;
                    16'h5FA2: data_out = 8'h3D;
                    16'h5FA3: data_out = 8'h3C;
                    16'h5FA4: data_out = 8'h3B;
                    16'h5FA5: data_out = 8'h3A;
                    16'h5FA6: data_out = 8'h39;
                    16'h5FA7: data_out = 8'h38;
                    16'h5FA8: data_out = 8'h37;
                    16'h5FA9: data_out = 8'h36;
                    16'h5FAA: data_out = 8'h35;
                    16'h5FAB: data_out = 8'h34;
                    16'h5FAC: data_out = 8'h33;
                    16'h5FAD: data_out = 8'h32;
                    16'h5FAE: data_out = 8'h31;
                    16'h5FAF: data_out = 8'h30;
                    16'h5FB0: data_out = 8'h2F;
                    16'h5FB1: data_out = 8'h2E;
                    16'h5FB2: data_out = 8'h2D;
                    16'h5FB3: data_out = 8'h2C;
                    16'h5FB4: data_out = 8'h2B;
                    16'h5FB5: data_out = 8'h2A;
                    16'h5FB6: data_out = 8'h29;
                    16'h5FB7: data_out = 8'h28;
                    16'h5FB8: data_out = 8'h27;
                    16'h5FB9: data_out = 8'h26;
                    16'h5FBA: data_out = 8'h25;
                    16'h5FBB: data_out = 8'h24;
                    16'h5FBC: data_out = 8'h23;
                    16'h5FBD: data_out = 8'h22;
                    16'h5FBE: data_out = 8'h21;
                    16'h5FBF: data_out = 8'h20;
                    16'h5FC0: data_out = 8'h1F;
                    16'h5FC1: data_out = 8'h1E;
                    16'h5FC2: data_out = 8'h1D;
                    16'h5FC3: data_out = 8'h1C;
                    16'h5FC4: data_out = 8'h1B;
                    16'h5FC5: data_out = 8'h1A;
                    16'h5FC6: data_out = 8'h19;
                    16'h5FC7: data_out = 8'h18;
                    16'h5FC8: data_out = 8'h17;
                    16'h5FC9: data_out = 8'h16;
                    16'h5FCA: data_out = 8'h15;
                    16'h5FCB: data_out = 8'h14;
                    16'h5FCC: data_out = 8'h13;
                    16'h5FCD: data_out = 8'h12;
                    16'h5FCE: data_out = 8'h11;
                    16'h5FCF: data_out = 8'h10;
                    16'h5FD0: data_out = 8'hF;
                    16'h5FD1: data_out = 8'hE;
                    16'h5FD2: data_out = 8'hD;
                    16'h5FD3: data_out = 8'hC;
                    16'h5FD4: data_out = 8'hB;
                    16'h5FD5: data_out = 8'hA;
                    16'h5FD6: data_out = 8'h9;
                    16'h5FD7: data_out = 8'h8;
                    16'h5FD8: data_out = 8'h7;
                    16'h5FD9: data_out = 8'h6;
                    16'h5FDA: data_out = 8'h5;
                    16'h5FDB: data_out = 8'h4;
                    16'h5FDC: data_out = 8'h3;
                    16'h5FDD: data_out = 8'h2;
                    16'h5FDE: data_out = 8'h1;
                    16'h5FDF: data_out = 8'h0;
                    16'h5FE0: data_out = 8'h81;
                    16'h5FE1: data_out = 8'h82;
                    16'h5FE2: data_out = 8'h83;
                    16'h5FE3: data_out = 8'h84;
                    16'h5FE4: data_out = 8'h85;
                    16'h5FE5: data_out = 8'h86;
                    16'h5FE6: data_out = 8'h87;
                    16'h5FE7: data_out = 8'h88;
                    16'h5FE8: data_out = 8'h89;
                    16'h5FE9: data_out = 8'h8A;
                    16'h5FEA: data_out = 8'h8B;
                    16'h5FEB: data_out = 8'h8C;
                    16'h5FEC: data_out = 8'h8D;
                    16'h5FED: data_out = 8'h8E;
                    16'h5FEE: data_out = 8'h8F;
                    16'h5FEF: data_out = 8'h90;
                    16'h5FF0: data_out = 8'h91;
                    16'h5FF1: data_out = 8'h92;
                    16'h5FF2: data_out = 8'h93;
                    16'h5FF3: data_out = 8'h94;
                    16'h5FF4: data_out = 8'h95;
                    16'h5FF5: data_out = 8'h96;
                    16'h5FF6: data_out = 8'h97;
                    16'h5FF7: data_out = 8'h98;
                    16'h5FF8: data_out = 8'h99;
                    16'h5FF9: data_out = 8'h9A;
                    16'h5FFA: data_out = 8'h9B;
                    16'h5FFB: data_out = 8'h9C;
                    16'h5FFC: data_out = 8'h9D;
                    16'h5FFD: data_out = 8'h9E;
                    16'h5FFE: data_out = 8'h9F;
                    16'h5FFF: data_out = 8'hA0;
                    16'h6000: data_out = 8'h60;
                    16'h6001: data_out = 8'h61;
                    16'h6002: data_out = 8'h62;
                    16'h6003: data_out = 8'h63;
                    16'h6004: data_out = 8'h64;
                    16'h6005: data_out = 8'h65;
                    16'h6006: data_out = 8'h66;
                    16'h6007: data_out = 8'h67;
                    16'h6008: data_out = 8'h68;
                    16'h6009: data_out = 8'h69;
                    16'h600A: data_out = 8'h6A;
                    16'h600B: data_out = 8'h6B;
                    16'h600C: data_out = 8'h6C;
                    16'h600D: data_out = 8'h6D;
                    16'h600E: data_out = 8'h6E;
                    16'h600F: data_out = 8'h6F;
                    16'h6010: data_out = 8'h70;
                    16'h6011: data_out = 8'h71;
                    16'h6012: data_out = 8'h72;
                    16'h6013: data_out = 8'h73;
                    16'h6014: data_out = 8'h74;
                    16'h6015: data_out = 8'h75;
                    16'h6016: data_out = 8'h76;
                    16'h6017: data_out = 8'h77;
                    16'h6018: data_out = 8'h78;
                    16'h6019: data_out = 8'h79;
                    16'h601A: data_out = 8'h7A;
                    16'h601B: data_out = 8'h7B;
                    16'h601C: data_out = 8'h7C;
                    16'h601D: data_out = 8'h7D;
                    16'h601E: data_out = 8'h7E;
                    16'h601F: data_out = 8'h7F;
                    16'h6020: data_out = 8'h80;
                    16'h6021: data_out = 8'h81;
                    16'h6022: data_out = 8'h82;
                    16'h6023: data_out = 8'h83;
                    16'h6024: data_out = 8'h84;
                    16'h6025: data_out = 8'h85;
                    16'h6026: data_out = 8'h86;
                    16'h6027: data_out = 8'h87;
                    16'h6028: data_out = 8'h88;
                    16'h6029: data_out = 8'h89;
                    16'h602A: data_out = 8'h8A;
                    16'h602B: data_out = 8'h8B;
                    16'h602C: data_out = 8'h8C;
                    16'h602D: data_out = 8'h8D;
                    16'h602E: data_out = 8'h8E;
                    16'h602F: data_out = 8'h8F;
                    16'h6030: data_out = 8'h90;
                    16'h6031: data_out = 8'h91;
                    16'h6032: data_out = 8'h92;
                    16'h6033: data_out = 8'h93;
                    16'h6034: data_out = 8'h94;
                    16'h6035: data_out = 8'h95;
                    16'h6036: data_out = 8'h96;
                    16'h6037: data_out = 8'h97;
                    16'h6038: data_out = 8'h98;
                    16'h6039: data_out = 8'h99;
                    16'h603A: data_out = 8'h9A;
                    16'h603B: data_out = 8'h9B;
                    16'h603C: data_out = 8'h9C;
                    16'h603D: data_out = 8'h9D;
                    16'h603E: data_out = 8'h9E;
                    16'h603F: data_out = 8'h9F;
                    16'h6040: data_out = 8'hA0;
                    16'h6041: data_out = 8'hA1;
                    16'h6042: data_out = 8'hA2;
                    16'h6043: data_out = 8'hA3;
                    16'h6044: data_out = 8'hA4;
                    16'h6045: data_out = 8'hA5;
                    16'h6046: data_out = 8'hA6;
                    16'h6047: data_out = 8'hA7;
                    16'h6048: data_out = 8'hA8;
                    16'h6049: data_out = 8'hA9;
                    16'h604A: data_out = 8'hAA;
                    16'h604B: data_out = 8'hAB;
                    16'h604C: data_out = 8'hAC;
                    16'h604D: data_out = 8'hAD;
                    16'h604E: data_out = 8'hAE;
                    16'h604F: data_out = 8'hAF;
                    16'h6050: data_out = 8'hB0;
                    16'h6051: data_out = 8'hB1;
                    16'h6052: data_out = 8'hB2;
                    16'h6053: data_out = 8'hB3;
                    16'h6054: data_out = 8'hB4;
                    16'h6055: data_out = 8'hB5;
                    16'h6056: data_out = 8'hB6;
                    16'h6057: data_out = 8'hB7;
                    16'h6058: data_out = 8'hB8;
                    16'h6059: data_out = 8'hB9;
                    16'h605A: data_out = 8'hBA;
                    16'h605B: data_out = 8'hBB;
                    16'h605C: data_out = 8'hBC;
                    16'h605D: data_out = 8'hBD;
                    16'h605E: data_out = 8'hBE;
                    16'h605F: data_out = 8'hBF;
                    16'h6060: data_out = 8'hC0;
                    16'h6061: data_out = 8'hC1;
                    16'h6062: data_out = 8'hC2;
                    16'h6063: data_out = 8'hC3;
                    16'h6064: data_out = 8'hC4;
                    16'h6065: data_out = 8'hC5;
                    16'h6066: data_out = 8'hC6;
                    16'h6067: data_out = 8'hC7;
                    16'h6068: data_out = 8'hC8;
                    16'h6069: data_out = 8'hC9;
                    16'h606A: data_out = 8'hCA;
                    16'h606B: data_out = 8'hCB;
                    16'h606C: data_out = 8'hCC;
                    16'h606D: data_out = 8'hCD;
                    16'h606E: data_out = 8'hCE;
                    16'h606F: data_out = 8'hCF;
                    16'h6070: data_out = 8'hD0;
                    16'h6071: data_out = 8'hD1;
                    16'h6072: data_out = 8'hD2;
                    16'h6073: data_out = 8'hD3;
                    16'h6074: data_out = 8'hD4;
                    16'h6075: data_out = 8'hD5;
                    16'h6076: data_out = 8'hD6;
                    16'h6077: data_out = 8'hD7;
                    16'h6078: data_out = 8'hD8;
                    16'h6079: data_out = 8'hD9;
                    16'h607A: data_out = 8'hDA;
                    16'h607B: data_out = 8'hDB;
                    16'h607C: data_out = 8'hDC;
                    16'h607D: data_out = 8'hDD;
                    16'h607E: data_out = 8'hDE;
                    16'h607F: data_out = 8'hDF;
                    16'h6080: data_out = 8'h60;
                    16'h6081: data_out = 8'h5F;
                    16'h6082: data_out = 8'h5E;
                    16'h6083: data_out = 8'h5D;
                    16'h6084: data_out = 8'h5C;
                    16'h6085: data_out = 8'h5B;
                    16'h6086: data_out = 8'h5A;
                    16'h6087: data_out = 8'h59;
                    16'h6088: data_out = 8'h58;
                    16'h6089: data_out = 8'h57;
                    16'h608A: data_out = 8'h56;
                    16'h608B: data_out = 8'h55;
                    16'h608C: data_out = 8'h54;
                    16'h608D: data_out = 8'h53;
                    16'h608E: data_out = 8'h52;
                    16'h608F: data_out = 8'h51;
                    16'h6090: data_out = 8'h50;
                    16'h6091: data_out = 8'h4F;
                    16'h6092: data_out = 8'h4E;
                    16'h6093: data_out = 8'h4D;
                    16'h6094: data_out = 8'h4C;
                    16'h6095: data_out = 8'h4B;
                    16'h6096: data_out = 8'h4A;
                    16'h6097: data_out = 8'h49;
                    16'h6098: data_out = 8'h48;
                    16'h6099: data_out = 8'h47;
                    16'h609A: data_out = 8'h46;
                    16'h609B: data_out = 8'h45;
                    16'h609C: data_out = 8'h44;
                    16'h609D: data_out = 8'h43;
                    16'h609E: data_out = 8'h42;
                    16'h609F: data_out = 8'h41;
                    16'h60A0: data_out = 8'h40;
                    16'h60A1: data_out = 8'h3F;
                    16'h60A2: data_out = 8'h3E;
                    16'h60A3: data_out = 8'h3D;
                    16'h60A4: data_out = 8'h3C;
                    16'h60A5: data_out = 8'h3B;
                    16'h60A6: data_out = 8'h3A;
                    16'h60A7: data_out = 8'h39;
                    16'h60A8: data_out = 8'h38;
                    16'h60A9: data_out = 8'h37;
                    16'h60AA: data_out = 8'h36;
                    16'h60AB: data_out = 8'h35;
                    16'h60AC: data_out = 8'h34;
                    16'h60AD: data_out = 8'h33;
                    16'h60AE: data_out = 8'h32;
                    16'h60AF: data_out = 8'h31;
                    16'h60B0: data_out = 8'h30;
                    16'h60B1: data_out = 8'h2F;
                    16'h60B2: data_out = 8'h2E;
                    16'h60B3: data_out = 8'h2D;
                    16'h60B4: data_out = 8'h2C;
                    16'h60B5: data_out = 8'h2B;
                    16'h60B6: data_out = 8'h2A;
                    16'h60B7: data_out = 8'h29;
                    16'h60B8: data_out = 8'h28;
                    16'h60B9: data_out = 8'h27;
                    16'h60BA: data_out = 8'h26;
                    16'h60BB: data_out = 8'h25;
                    16'h60BC: data_out = 8'h24;
                    16'h60BD: data_out = 8'h23;
                    16'h60BE: data_out = 8'h22;
                    16'h60BF: data_out = 8'h21;
                    16'h60C0: data_out = 8'h20;
                    16'h60C1: data_out = 8'h1F;
                    16'h60C2: data_out = 8'h1E;
                    16'h60C3: data_out = 8'h1D;
                    16'h60C4: data_out = 8'h1C;
                    16'h60C5: data_out = 8'h1B;
                    16'h60C6: data_out = 8'h1A;
                    16'h60C7: data_out = 8'h19;
                    16'h60C8: data_out = 8'h18;
                    16'h60C9: data_out = 8'h17;
                    16'h60CA: data_out = 8'h16;
                    16'h60CB: data_out = 8'h15;
                    16'h60CC: data_out = 8'h14;
                    16'h60CD: data_out = 8'h13;
                    16'h60CE: data_out = 8'h12;
                    16'h60CF: data_out = 8'h11;
                    16'h60D0: data_out = 8'h10;
                    16'h60D1: data_out = 8'hF;
                    16'h60D2: data_out = 8'hE;
                    16'h60D3: data_out = 8'hD;
                    16'h60D4: data_out = 8'hC;
                    16'h60D5: data_out = 8'hB;
                    16'h60D6: data_out = 8'hA;
                    16'h60D7: data_out = 8'h9;
                    16'h60D8: data_out = 8'h8;
                    16'h60D9: data_out = 8'h7;
                    16'h60DA: data_out = 8'h6;
                    16'h60DB: data_out = 8'h5;
                    16'h60DC: data_out = 8'h4;
                    16'h60DD: data_out = 8'h3;
                    16'h60DE: data_out = 8'h2;
                    16'h60DF: data_out = 8'h1;
                    16'h60E0: data_out = 8'h0;
                    16'h60E1: data_out = 8'h81;
                    16'h60E2: data_out = 8'h82;
                    16'h60E3: data_out = 8'h83;
                    16'h60E4: data_out = 8'h84;
                    16'h60E5: data_out = 8'h85;
                    16'h60E6: data_out = 8'h86;
                    16'h60E7: data_out = 8'h87;
                    16'h60E8: data_out = 8'h88;
                    16'h60E9: data_out = 8'h89;
                    16'h60EA: data_out = 8'h8A;
                    16'h60EB: data_out = 8'h8B;
                    16'h60EC: data_out = 8'h8C;
                    16'h60ED: data_out = 8'h8D;
                    16'h60EE: data_out = 8'h8E;
                    16'h60EF: data_out = 8'h8F;
                    16'h60F0: data_out = 8'h90;
                    16'h60F1: data_out = 8'h91;
                    16'h60F2: data_out = 8'h92;
                    16'h60F3: data_out = 8'h93;
                    16'h60F4: data_out = 8'h94;
                    16'h60F5: data_out = 8'h95;
                    16'h60F6: data_out = 8'h96;
                    16'h60F7: data_out = 8'h97;
                    16'h60F8: data_out = 8'h98;
                    16'h60F9: data_out = 8'h99;
                    16'h60FA: data_out = 8'h9A;
                    16'h60FB: data_out = 8'h9B;
                    16'h60FC: data_out = 8'h9C;
                    16'h60FD: data_out = 8'h9D;
                    16'h60FE: data_out = 8'h9E;
                    16'h60FF: data_out = 8'h9F;
                    16'h6100: data_out = 8'h61;
                    16'h6101: data_out = 8'h62;
                    16'h6102: data_out = 8'h63;
                    16'h6103: data_out = 8'h64;
                    16'h6104: data_out = 8'h65;
                    16'h6105: data_out = 8'h66;
                    16'h6106: data_out = 8'h67;
                    16'h6107: data_out = 8'h68;
                    16'h6108: data_out = 8'h69;
                    16'h6109: data_out = 8'h6A;
                    16'h610A: data_out = 8'h6B;
                    16'h610B: data_out = 8'h6C;
                    16'h610C: data_out = 8'h6D;
                    16'h610D: data_out = 8'h6E;
                    16'h610E: data_out = 8'h6F;
                    16'h610F: data_out = 8'h70;
                    16'h6110: data_out = 8'h71;
                    16'h6111: data_out = 8'h72;
                    16'h6112: data_out = 8'h73;
                    16'h6113: data_out = 8'h74;
                    16'h6114: data_out = 8'h75;
                    16'h6115: data_out = 8'h76;
                    16'h6116: data_out = 8'h77;
                    16'h6117: data_out = 8'h78;
                    16'h6118: data_out = 8'h79;
                    16'h6119: data_out = 8'h7A;
                    16'h611A: data_out = 8'h7B;
                    16'h611B: data_out = 8'h7C;
                    16'h611C: data_out = 8'h7D;
                    16'h611D: data_out = 8'h7E;
                    16'h611E: data_out = 8'h7F;
                    16'h611F: data_out = 8'h80;
                    16'h6120: data_out = 8'h81;
                    16'h6121: data_out = 8'h82;
                    16'h6122: data_out = 8'h83;
                    16'h6123: data_out = 8'h84;
                    16'h6124: data_out = 8'h85;
                    16'h6125: data_out = 8'h86;
                    16'h6126: data_out = 8'h87;
                    16'h6127: data_out = 8'h88;
                    16'h6128: data_out = 8'h89;
                    16'h6129: data_out = 8'h8A;
                    16'h612A: data_out = 8'h8B;
                    16'h612B: data_out = 8'h8C;
                    16'h612C: data_out = 8'h8D;
                    16'h612D: data_out = 8'h8E;
                    16'h612E: data_out = 8'h8F;
                    16'h612F: data_out = 8'h90;
                    16'h6130: data_out = 8'h91;
                    16'h6131: data_out = 8'h92;
                    16'h6132: data_out = 8'h93;
                    16'h6133: data_out = 8'h94;
                    16'h6134: data_out = 8'h95;
                    16'h6135: data_out = 8'h96;
                    16'h6136: data_out = 8'h97;
                    16'h6137: data_out = 8'h98;
                    16'h6138: data_out = 8'h99;
                    16'h6139: data_out = 8'h9A;
                    16'h613A: data_out = 8'h9B;
                    16'h613B: data_out = 8'h9C;
                    16'h613C: data_out = 8'h9D;
                    16'h613D: data_out = 8'h9E;
                    16'h613E: data_out = 8'h9F;
                    16'h613F: data_out = 8'hA0;
                    16'h6140: data_out = 8'hA1;
                    16'h6141: data_out = 8'hA2;
                    16'h6142: data_out = 8'hA3;
                    16'h6143: data_out = 8'hA4;
                    16'h6144: data_out = 8'hA5;
                    16'h6145: data_out = 8'hA6;
                    16'h6146: data_out = 8'hA7;
                    16'h6147: data_out = 8'hA8;
                    16'h6148: data_out = 8'hA9;
                    16'h6149: data_out = 8'hAA;
                    16'h614A: data_out = 8'hAB;
                    16'h614B: data_out = 8'hAC;
                    16'h614C: data_out = 8'hAD;
                    16'h614D: data_out = 8'hAE;
                    16'h614E: data_out = 8'hAF;
                    16'h614F: data_out = 8'hB0;
                    16'h6150: data_out = 8'hB1;
                    16'h6151: data_out = 8'hB2;
                    16'h6152: data_out = 8'hB3;
                    16'h6153: data_out = 8'hB4;
                    16'h6154: data_out = 8'hB5;
                    16'h6155: data_out = 8'hB6;
                    16'h6156: data_out = 8'hB7;
                    16'h6157: data_out = 8'hB8;
                    16'h6158: data_out = 8'hB9;
                    16'h6159: data_out = 8'hBA;
                    16'h615A: data_out = 8'hBB;
                    16'h615B: data_out = 8'hBC;
                    16'h615C: data_out = 8'hBD;
                    16'h615D: data_out = 8'hBE;
                    16'h615E: data_out = 8'hBF;
                    16'h615F: data_out = 8'hC0;
                    16'h6160: data_out = 8'hC1;
                    16'h6161: data_out = 8'hC2;
                    16'h6162: data_out = 8'hC3;
                    16'h6163: data_out = 8'hC4;
                    16'h6164: data_out = 8'hC5;
                    16'h6165: data_out = 8'hC6;
                    16'h6166: data_out = 8'hC7;
                    16'h6167: data_out = 8'hC8;
                    16'h6168: data_out = 8'hC9;
                    16'h6169: data_out = 8'hCA;
                    16'h616A: data_out = 8'hCB;
                    16'h616B: data_out = 8'hCC;
                    16'h616C: data_out = 8'hCD;
                    16'h616D: data_out = 8'hCE;
                    16'h616E: data_out = 8'hCF;
                    16'h616F: data_out = 8'hD0;
                    16'h6170: data_out = 8'hD1;
                    16'h6171: data_out = 8'hD2;
                    16'h6172: data_out = 8'hD3;
                    16'h6173: data_out = 8'hD4;
                    16'h6174: data_out = 8'hD5;
                    16'h6175: data_out = 8'hD6;
                    16'h6176: data_out = 8'hD7;
                    16'h6177: data_out = 8'hD8;
                    16'h6178: data_out = 8'hD9;
                    16'h6179: data_out = 8'hDA;
                    16'h617A: data_out = 8'hDB;
                    16'h617B: data_out = 8'hDC;
                    16'h617C: data_out = 8'hDD;
                    16'h617D: data_out = 8'hDE;
                    16'h617E: data_out = 8'hDF;
                    16'h617F: data_out = 8'hE0;
                    16'h6180: data_out = 8'h61;
                    16'h6181: data_out = 8'h60;
                    16'h6182: data_out = 8'h5F;
                    16'h6183: data_out = 8'h5E;
                    16'h6184: data_out = 8'h5D;
                    16'h6185: data_out = 8'h5C;
                    16'h6186: data_out = 8'h5B;
                    16'h6187: data_out = 8'h5A;
                    16'h6188: data_out = 8'h59;
                    16'h6189: data_out = 8'h58;
                    16'h618A: data_out = 8'h57;
                    16'h618B: data_out = 8'h56;
                    16'h618C: data_out = 8'h55;
                    16'h618D: data_out = 8'h54;
                    16'h618E: data_out = 8'h53;
                    16'h618F: data_out = 8'h52;
                    16'h6190: data_out = 8'h51;
                    16'h6191: data_out = 8'h50;
                    16'h6192: data_out = 8'h4F;
                    16'h6193: data_out = 8'h4E;
                    16'h6194: data_out = 8'h4D;
                    16'h6195: data_out = 8'h4C;
                    16'h6196: data_out = 8'h4B;
                    16'h6197: data_out = 8'h4A;
                    16'h6198: data_out = 8'h49;
                    16'h6199: data_out = 8'h48;
                    16'h619A: data_out = 8'h47;
                    16'h619B: data_out = 8'h46;
                    16'h619C: data_out = 8'h45;
                    16'h619D: data_out = 8'h44;
                    16'h619E: data_out = 8'h43;
                    16'h619F: data_out = 8'h42;
                    16'h61A0: data_out = 8'h41;
                    16'h61A1: data_out = 8'h40;
                    16'h61A2: data_out = 8'h3F;
                    16'h61A3: data_out = 8'h3E;
                    16'h61A4: data_out = 8'h3D;
                    16'h61A5: data_out = 8'h3C;
                    16'h61A6: data_out = 8'h3B;
                    16'h61A7: data_out = 8'h3A;
                    16'h61A8: data_out = 8'h39;
                    16'h61A9: data_out = 8'h38;
                    16'h61AA: data_out = 8'h37;
                    16'h61AB: data_out = 8'h36;
                    16'h61AC: data_out = 8'h35;
                    16'h61AD: data_out = 8'h34;
                    16'h61AE: data_out = 8'h33;
                    16'h61AF: data_out = 8'h32;
                    16'h61B0: data_out = 8'h31;
                    16'h61B1: data_out = 8'h30;
                    16'h61B2: data_out = 8'h2F;
                    16'h61B3: data_out = 8'h2E;
                    16'h61B4: data_out = 8'h2D;
                    16'h61B5: data_out = 8'h2C;
                    16'h61B6: data_out = 8'h2B;
                    16'h61B7: data_out = 8'h2A;
                    16'h61B8: data_out = 8'h29;
                    16'h61B9: data_out = 8'h28;
                    16'h61BA: data_out = 8'h27;
                    16'h61BB: data_out = 8'h26;
                    16'h61BC: data_out = 8'h25;
                    16'h61BD: data_out = 8'h24;
                    16'h61BE: data_out = 8'h23;
                    16'h61BF: data_out = 8'h22;
                    16'h61C0: data_out = 8'h21;
                    16'h61C1: data_out = 8'h20;
                    16'h61C2: data_out = 8'h1F;
                    16'h61C3: data_out = 8'h1E;
                    16'h61C4: data_out = 8'h1D;
                    16'h61C5: data_out = 8'h1C;
                    16'h61C6: data_out = 8'h1B;
                    16'h61C7: data_out = 8'h1A;
                    16'h61C8: data_out = 8'h19;
                    16'h61C9: data_out = 8'h18;
                    16'h61CA: data_out = 8'h17;
                    16'h61CB: data_out = 8'h16;
                    16'h61CC: data_out = 8'h15;
                    16'h61CD: data_out = 8'h14;
                    16'h61CE: data_out = 8'h13;
                    16'h61CF: data_out = 8'h12;
                    16'h61D0: data_out = 8'h11;
                    16'h61D1: data_out = 8'h10;
                    16'h61D2: data_out = 8'hF;
                    16'h61D3: data_out = 8'hE;
                    16'h61D4: data_out = 8'hD;
                    16'h61D5: data_out = 8'hC;
                    16'h61D6: data_out = 8'hB;
                    16'h61D7: data_out = 8'hA;
                    16'h61D8: data_out = 8'h9;
                    16'h61D9: data_out = 8'h8;
                    16'h61DA: data_out = 8'h7;
                    16'h61DB: data_out = 8'h6;
                    16'h61DC: data_out = 8'h5;
                    16'h61DD: data_out = 8'h4;
                    16'h61DE: data_out = 8'h3;
                    16'h61DF: data_out = 8'h2;
                    16'h61E0: data_out = 8'h1;
                    16'h61E1: data_out = 8'h0;
                    16'h61E2: data_out = 8'h81;
                    16'h61E3: data_out = 8'h82;
                    16'h61E4: data_out = 8'h83;
                    16'h61E5: data_out = 8'h84;
                    16'h61E6: data_out = 8'h85;
                    16'h61E7: data_out = 8'h86;
                    16'h61E8: data_out = 8'h87;
                    16'h61E9: data_out = 8'h88;
                    16'h61EA: data_out = 8'h89;
                    16'h61EB: data_out = 8'h8A;
                    16'h61EC: data_out = 8'h8B;
                    16'h61ED: data_out = 8'h8C;
                    16'h61EE: data_out = 8'h8D;
                    16'h61EF: data_out = 8'h8E;
                    16'h61F0: data_out = 8'h8F;
                    16'h61F1: data_out = 8'h90;
                    16'h61F2: data_out = 8'h91;
                    16'h61F3: data_out = 8'h92;
                    16'h61F4: data_out = 8'h93;
                    16'h61F5: data_out = 8'h94;
                    16'h61F6: data_out = 8'h95;
                    16'h61F7: data_out = 8'h96;
                    16'h61F8: data_out = 8'h97;
                    16'h61F9: data_out = 8'h98;
                    16'h61FA: data_out = 8'h99;
                    16'h61FB: data_out = 8'h9A;
                    16'h61FC: data_out = 8'h9B;
                    16'h61FD: data_out = 8'h9C;
                    16'h61FE: data_out = 8'h9D;
                    16'h61FF: data_out = 8'h9E;
                    16'h6200: data_out = 8'h62;
                    16'h6201: data_out = 8'h63;
                    16'h6202: data_out = 8'h64;
                    16'h6203: data_out = 8'h65;
                    16'h6204: data_out = 8'h66;
                    16'h6205: data_out = 8'h67;
                    16'h6206: data_out = 8'h68;
                    16'h6207: data_out = 8'h69;
                    16'h6208: data_out = 8'h6A;
                    16'h6209: data_out = 8'h6B;
                    16'h620A: data_out = 8'h6C;
                    16'h620B: data_out = 8'h6D;
                    16'h620C: data_out = 8'h6E;
                    16'h620D: data_out = 8'h6F;
                    16'h620E: data_out = 8'h70;
                    16'h620F: data_out = 8'h71;
                    16'h6210: data_out = 8'h72;
                    16'h6211: data_out = 8'h73;
                    16'h6212: data_out = 8'h74;
                    16'h6213: data_out = 8'h75;
                    16'h6214: data_out = 8'h76;
                    16'h6215: data_out = 8'h77;
                    16'h6216: data_out = 8'h78;
                    16'h6217: data_out = 8'h79;
                    16'h6218: data_out = 8'h7A;
                    16'h6219: data_out = 8'h7B;
                    16'h621A: data_out = 8'h7C;
                    16'h621B: data_out = 8'h7D;
                    16'h621C: data_out = 8'h7E;
                    16'h621D: data_out = 8'h7F;
                    16'h621E: data_out = 8'h80;
                    16'h621F: data_out = 8'h81;
                    16'h6220: data_out = 8'h82;
                    16'h6221: data_out = 8'h83;
                    16'h6222: data_out = 8'h84;
                    16'h6223: data_out = 8'h85;
                    16'h6224: data_out = 8'h86;
                    16'h6225: data_out = 8'h87;
                    16'h6226: data_out = 8'h88;
                    16'h6227: data_out = 8'h89;
                    16'h6228: data_out = 8'h8A;
                    16'h6229: data_out = 8'h8B;
                    16'h622A: data_out = 8'h8C;
                    16'h622B: data_out = 8'h8D;
                    16'h622C: data_out = 8'h8E;
                    16'h622D: data_out = 8'h8F;
                    16'h622E: data_out = 8'h90;
                    16'h622F: data_out = 8'h91;
                    16'h6230: data_out = 8'h92;
                    16'h6231: data_out = 8'h93;
                    16'h6232: data_out = 8'h94;
                    16'h6233: data_out = 8'h95;
                    16'h6234: data_out = 8'h96;
                    16'h6235: data_out = 8'h97;
                    16'h6236: data_out = 8'h98;
                    16'h6237: data_out = 8'h99;
                    16'h6238: data_out = 8'h9A;
                    16'h6239: data_out = 8'h9B;
                    16'h623A: data_out = 8'h9C;
                    16'h623B: data_out = 8'h9D;
                    16'h623C: data_out = 8'h9E;
                    16'h623D: data_out = 8'h9F;
                    16'h623E: data_out = 8'hA0;
                    16'h623F: data_out = 8'hA1;
                    16'h6240: data_out = 8'hA2;
                    16'h6241: data_out = 8'hA3;
                    16'h6242: data_out = 8'hA4;
                    16'h6243: data_out = 8'hA5;
                    16'h6244: data_out = 8'hA6;
                    16'h6245: data_out = 8'hA7;
                    16'h6246: data_out = 8'hA8;
                    16'h6247: data_out = 8'hA9;
                    16'h6248: data_out = 8'hAA;
                    16'h6249: data_out = 8'hAB;
                    16'h624A: data_out = 8'hAC;
                    16'h624B: data_out = 8'hAD;
                    16'h624C: data_out = 8'hAE;
                    16'h624D: data_out = 8'hAF;
                    16'h624E: data_out = 8'hB0;
                    16'h624F: data_out = 8'hB1;
                    16'h6250: data_out = 8'hB2;
                    16'h6251: data_out = 8'hB3;
                    16'h6252: data_out = 8'hB4;
                    16'h6253: data_out = 8'hB5;
                    16'h6254: data_out = 8'hB6;
                    16'h6255: data_out = 8'hB7;
                    16'h6256: data_out = 8'hB8;
                    16'h6257: data_out = 8'hB9;
                    16'h6258: data_out = 8'hBA;
                    16'h6259: data_out = 8'hBB;
                    16'h625A: data_out = 8'hBC;
                    16'h625B: data_out = 8'hBD;
                    16'h625C: data_out = 8'hBE;
                    16'h625D: data_out = 8'hBF;
                    16'h625E: data_out = 8'hC0;
                    16'h625F: data_out = 8'hC1;
                    16'h6260: data_out = 8'hC2;
                    16'h6261: data_out = 8'hC3;
                    16'h6262: data_out = 8'hC4;
                    16'h6263: data_out = 8'hC5;
                    16'h6264: data_out = 8'hC6;
                    16'h6265: data_out = 8'hC7;
                    16'h6266: data_out = 8'hC8;
                    16'h6267: data_out = 8'hC9;
                    16'h6268: data_out = 8'hCA;
                    16'h6269: data_out = 8'hCB;
                    16'h626A: data_out = 8'hCC;
                    16'h626B: data_out = 8'hCD;
                    16'h626C: data_out = 8'hCE;
                    16'h626D: data_out = 8'hCF;
                    16'h626E: data_out = 8'hD0;
                    16'h626F: data_out = 8'hD1;
                    16'h6270: data_out = 8'hD2;
                    16'h6271: data_out = 8'hD3;
                    16'h6272: data_out = 8'hD4;
                    16'h6273: data_out = 8'hD5;
                    16'h6274: data_out = 8'hD6;
                    16'h6275: data_out = 8'hD7;
                    16'h6276: data_out = 8'hD8;
                    16'h6277: data_out = 8'hD9;
                    16'h6278: data_out = 8'hDA;
                    16'h6279: data_out = 8'hDB;
                    16'h627A: data_out = 8'hDC;
                    16'h627B: data_out = 8'hDD;
                    16'h627C: data_out = 8'hDE;
                    16'h627D: data_out = 8'hDF;
                    16'h627E: data_out = 8'hE0;
                    16'h627F: data_out = 8'hE1;
                    16'h6280: data_out = 8'h62;
                    16'h6281: data_out = 8'h61;
                    16'h6282: data_out = 8'h60;
                    16'h6283: data_out = 8'h5F;
                    16'h6284: data_out = 8'h5E;
                    16'h6285: data_out = 8'h5D;
                    16'h6286: data_out = 8'h5C;
                    16'h6287: data_out = 8'h5B;
                    16'h6288: data_out = 8'h5A;
                    16'h6289: data_out = 8'h59;
                    16'h628A: data_out = 8'h58;
                    16'h628B: data_out = 8'h57;
                    16'h628C: data_out = 8'h56;
                    16'h628D: data_out = 8'h55;
                    16'h628E: data_out = 8'h54;
                    16'h628F: data_out = 8'h53;
                    16'h6290: data_out = 8'h52;
                    16'h6291: data_out = 8'h51;
                    16'h6292: data_out = 8'h50;
                    16'h6293: data_out = 8'h4F;
                    16'h6294: data_out = 8'h4E;
                    16'h6295: data_out = 8'h4D;
                    16'h6296: data_out = 8'h4C;
                    16'h6297: data_out = 8'h4B;
                    16'h6298: data_out = 8'h4A;
                    16'h6299: data_out = 8'h49;
                    16'h629A: data_out = 8'h48;
                    16'h629B: data_out = 8'h47;
                    16'h629C: data_out = 8'h46;
                    16'h629D: data_out = 8'h45;
                    16'h629E: data_out = 8'h44;
                    16'h629F: data_out = 8'h43;
                    16'h62A0: data_out = 8'h42;
                    16'h62A1: data_out = 8'h41;
                    16'h62A2: data_out = 8'h40;
                    16'h62A3: data_out = 8'h3F;
                    16'h62A4: data_out = 8'h3E;
                    16'h62A5: data_out = 8'h3D;
                    16'h62A6: data_out = 8'h3C;
                    16'h62A7: data_out = 8'h3B;
                    16'h62A8: data_out = 8'h3A;
                    16'h62A9: data_out = 8'h39;
                    16'h62AA: data_out = 8'h38;
                    16'h62AB: data_out = 8'h37;
                    16'h62AC: data_out = 8'h36;
                    16'h62AD: data_out = 8'h35;
                    16'h62AE: data_out = 8'h34;
                    16'h62AF: data_out = 8'h33;
                    16'h62B0: data_out = 8'h32;
                    16'h62B1: data_out = 8'h31;
                    16'h62B2: data_out = 8'h30;
                    16'h62B3: data_out = 8'h2F;
                    16'h62B4: data_out = 8'h2E;
                    16'h62B5: data_out = 8'h2D;
                    16'h62B6: data_out = 8'h2C;
                    16'h62B7: data_out = 8'h2B;
                    16'h62B8: data_out = 8'h2A;
                    16'h62B9: data_out = 8'h29;
                    16'h62BA: data_out = 8'h28;
                    16'h62BB: data_out = 8'h27;
                    16'h62BC: data_out = 8'h26;
                    16'h62BD: data_out = 8'h25;
                    16'h62BE: data_out = 8'h24;
                    16'h62BF: data_out = 8'h23;
                    16'h62C0: data_out = 8'h22;
                    16'h62C1: data_out = 8'h21;
                    16'h62C2: data_out = 8'h20;
                    16'h62C3: data_out = 8'h1F;
                    16'h62C4: data_out = 8'h1E;
                    16'h62C5: data_out = 8'h1D;
                    16'h62C6: data_out = 8'h1C;
                    16'h62C7: data_out = 8'h1B;
                    16'h62C8: data_out = 8'h1A;
                    16'h62C9: data_out = 8'h19;
                    16'h62CA: data_out = 8'h18;
                    16'h62CB: data_out = 8'h17;
                    16'h62CC: data_out = 8'h16;
                    16'h62CD: data_out = 8'h15;
                    16'h62CE: data_out = 8'h14;
                    16'h62CF: data_out = 8'h13;
                    16'h62D0: data_out = 8'h12;
                    16'h62D1: data_out = 8'h11;
                    16'h62D2: data_out = 8'h10;
                    16'h62D3: data_out = 8'hF;
                    16'h62D4: data_out = 8'hE;
                    16'h62D5: data_out = 8'hD;
                    16'h62D6: data_out = 8'hC;
                    16'h62D7: data_out = 8'hB;
                    16'h62D8: data_out = 8'hA;
                    16'h62D9: data_out = 8'h9;
                    16'h62DA: data_out = 8'h8;
                    16'h62DB: data_out = 8'h7;
                    16'h62DC: data_out = 8'h6;
                    16'h62DD: data_out = 8'h5;
                    16'h62DE: data_out = 8'h4;
                    16'h62DF: data_out = 8'h3;
                    16'h62E0: data_out = 8'h2;
                    16'h62E1: data_out = 8'h1;
                    16'h62E2: data_out = 8'h0;
                    16'h62E3: data_out = 8'h81;
                    16'h62E4: data_out = 8'h82;
                    16'h62E5: data_out = 8'h83;
                    16'h62E6: data_out = 8'h84;
                    16'h62E7: data_out = 8'h85;
                    16'h62E8: data_out = 8'h86;
                    16'h62E9: data_out = 8'h87;
                    16'h62EA: data_out = 8'h88;
                    16'h62EB: data_out = 8'h89;
                    16'h62EC: data_out = 8'h8A;
                    16'h62ED: data_out = 8'h8B;
                    16'h62EE: data_out = 8'h8C;
                    16'h62EF: data_out = 8'h8D;
                    16'h62F0: data_out = 8'h8E;
                    16'h62F1: data_out = 8'h8F;
                    16'h62F2: data_out = 8'h90;
                    16'h62F3: data_out = 8'h91;
                    16'h62F4: data_out = 8'h92;
                    16'h62F5: data_out = 8'h93;
                    16'h62F6: data_out = 8'h94;
                    16'h62F7: data_out = 8'h95;
                    16'h62F8: data_out = 8'h96;
                    16'h62F9: data_out = 8'h97;
                    16'h62FA: data_out = 8'h98;
                    16'h62FB: data_out = 8'h99;
                    16'h62FC: data_out = 8'h9A;
                    16'h62FD: data_out = 8'h9B;
                    16'h62FE: data_out = 8'h9C;
                    16'h62FF: data_out = 8'h9D;
                    16'h6300: data_out = 8'h63;
                    16'h6301: data_out = 8'h64;
                    16'h6302: data_out = 8'h65;
                    16'h6303: data_out = 8'h66;
                    16'h6304: data_out = 8'h67;
                    16'h6305: data_out = 8'h68;
                    16'h6306: data_out = 8'h69;
                    16'h6307: data_out = 8'h6A;
                    16'h6308: data_out = 8'h6B;
                    16'h6309: data_out = 8'h6C;
                    16'h630A: data_out = 8'h6D;
                    16'h630B: data_out = 8'h6E;
                    16'h630C: data_out = 8'h6F;
                    16'h630D: data_out = 8'h70;
                    16'h630E: data_out = 8'h71;
                    16'h630F: data_out = 8'h72;
                    16'h6310: data_out = 8'h73;
                    16'h6311: data_out = 8'h74;
                    16'h6312: data_out = 8'h75;
                    16'h6313: data_out = 8'h76;
                    16'h6314: data_out = 8'h77;
                    16'h6315: data_out = 8'h78;
                    16'h6316: data_out = 8'h79;
                    16'h6317: data_out = 8'h7A;
                    16'h6318: data_out = 8'h7B;
                    16'h6319: data_out = 8'h7C;
                    16'h631A: data_out = 8'h7D;
                    16'h631B: data_out = 8'h7E;
                    16'h631C: data_out = 8'h7F;
                    16'h631D: data_out = 8'h80;
                    16'h631E: data_out = 8'h81;
                    16'h631F: data_out = 8'h82;
                    16'h6320: data_out = 8'h83;
                    16'h6321: data_out = 8'h84;
                    16'h6322: data_out = 8'h85;
                    16'h6323: data_out = 8'h86;
                    16'h6324: data_out = 8'h87;
                    16'h6325: data_out = 8'h88;
                    16'h6326: data_out = 8'h89;
                    16'h6327: data_out = 8'h8A;
                    16'h6328: data_out = 8'h8B;
                    16'h6329: data_out = 8'h8C;
                    16'h632A: data_out = 8'h8D;
                    16'h632B: data_out = 8'h8E;
                    16'h632C: data_out = 8'h8F;
                    16'h632D: data_out = 8'h90;
                    16'h632E: data_out = 8'h91;
                    16'h632F: data_out = 8'h92;
                    16'h6330: data_out = 8'h93;
                    16'h6331: data_out = 8'h94;
                    16'h6332: data_out = 8'h95;
                    16'h6333: data_out = 8'h96;
                    16'h6334: data_out = 8'h97;
                    16'h6335: data_out = 8'h98;
                    16'h6336: data_out = 8'h99;
                    16'h6337: data_out = 8'h9A;
                    16'h6338: data_out = 8'h9B;
                    16'h6339: data_out = 8'h9C;
                    16'h633A: data_out = 8'h9D;
                    16'h633B: data_out = 8'h9E;
                    16'h633C: data_out = 8'h9F;
                    16'h633D: data_out = 8'hA0;
                    16'h633E: data_out = 8'hA1;
                    16'h633F: data_out = 8'hA2;
                    16'h6340: data_out = 8'hA3;
                    16'h6341: data_out = 8'hA4;
                    16'h6342: data_out = 8'hA5;
                    16'h6343: data_out = 8'hA6;
                    16'h6344: data_out = 8'hA7;
                    16'h6345: data_out = 8'hA8;
                    16'h6346: data_out = 8'hA9;
                    16'h6347: data_out = 8'hAA;
                    16'h6348: data_out = 8'hAB;
                    16'h6349: data_out = 8'hAC;
                    16'h634A: data_out = 8'hAD;
                    16'h634B: data_out = 8'hAE;
                    16'h634C: data_out = 8'hAF;
                    16'h634D: data_out = 8'hB0;
                    16'h634E: data_out = 8'hB1;
                    16'h634F: data_out = 8'hB2;
                    16'h6350: data_out = 8'hB3;
                    16'h6351: data_out = 8'hB4;
                    16'h6352: data_out = 8'hB5;
                    16'h6353: data_out = 8'hB6;
                    16'h6354: data_out = 8'hB7;
                    16'h6355: data_out = 8'hB8;
                    16'h6356: data_out = 8'hB9;
                    16'h6357: data_out = 8'hBA;
                    16'h6358: data_out = 8'hBB;
                    16'h6359: data_out = 8'hBC;
                    16'h635A: data_out = 8'hBD;
                    16'h635B: data_out = 8'hBE;
                    16'h635C: data_out = 8'hBF;
                    16'h635D: data_out = 8'hC0;
                    16'h635E: data_out = 8'hC1;
                    16'h635F: data_out = 8'hC2;
                    16'h6360: data_out = 8'hC3;
                    16'h6361: data_out = 8'hC4;
                    16'h6362: data_out = 8'hC5;
                    16'h6363: data_out = 8'hC6;
                    16'h6364: data_out = 8'hC7;
                    16'h6365: data_out = 8'hC8;
                    16'h6366: data_out = 8'hC9;
                    16'h6367: data_out = 8'hCA;
                    16'h6368: data_out = 8'hCB;
                    16'h6369: data_out = 8'hCC;
                    16'h636A: data_out = 8'hCD;
                    16'h636B: data_out = 8'hCE;
                    16'h636C: data_out = 8'hCF;
                    16'h636D: data_out = 8'hD0;
                    16'h636E: data_out = 8'hD1;
                    16'h636F: data_out = 8'hD2;
                    16'h6370: data_out = 8'hD3;
                    16'h6371: data_out = 8'hD4;
                    16'h6372: data_out = 8'hD5;
                    16'h6373: data_out = 8'hD6;
                    16'h6374: data_out = 8'hD7;
                    16'h6375: data_out = 8'hD8;
                    16'h6376: data_out = 8'hD9;
                    16'h6377: data_out = 8'hDA;
                    16'h6378: data_out = 8'hDB;
                    16'h6379: data_out = 8'hDC;
                    16'h637A: data_out = 8'hDD;
                    16'h637B: data_out = 8'hDE;
                    16'h637C: data_out = 8'hDF;
                    16'h637D: data_out = 8'hE0;
                    16'h637E: data_out = 8'hE1;
                    16'h637F: data_out = 8'hE2;
                    16'h6380: data_out = 8'h63;
                    16'h6381: data_out = 8'h62;
                    16'h6382: data_out = 8'h61;
                    16'h6383: data_out = 8'h60;
                    16'h6384: data_out = 8'h5F;
                    16'h6385: data_out = 8'h5E;
                    16'h6386: data_out = 8'h5D;
                    16'h6387: data_out = 8'h5C;
                    16'h6388: data_out = 8'h5B;
                    16'h6389: data_out = 8'h5A;
                    16'h638A: data_out = 8'h59;
                    16'h638B: data_out = 8'h58;
                    16'h638C: data_out = 8'h57;
                    16'h638D: data_out = 8'h56;
                    16'h638E: data_out = 8'h55;
                    16'h638F: data_out = 8'h54;
                    16'h6390: data_out = 8'h53;
                    16'h6391: data_out = 8'h52;
                    16'h6392: data_out = 8'h51;
                    16'h6393: data_out = 8'h50;
                    16'h6394: data_out = 8'h4F;
                    16'h6395: data_out = 8'h4E;
                    16'h6396: data_out = 8'h4D;
                    16'h6397: data_out = 8'h4C;
                    16'h6398: data_out = 8'h4B;
                    16'h6399: data_out = 8'h4A;
                    16'h639A: data_out = 8'h49;
                    16'h639B: data_out = 8'h48;
                    16'h639C: data_out = 8'h47;
                    16'h639D: data_out = 8'h46;
                    16'h639E: data_out = 8'h45;
                    16'h639F: data_out = 8'h44;
                    16'h63A0: data_out = 8'h43;
                    16'h63A1: data_out = 8'h42;
                    16'h63A2: data_out = 8'h41;
                    16'h63A3: data_out = 8'h40;
                    16'h63A4: data_out = 8'h3F;
                    16'h63A5: data_out = 8'h3E;
                    16'h63A6: data_out = 8'h3D;
                    16'h63A7: data_out = 8'h3C;
                    16'h63A8: data_out = 8'h3B;
                    16'h63A9: data_out = 8'h3A;
                    16'h63AA: data_out = 8'h39;
                    16'h63AB: data_out = 8'h38;
                    16'h63AC: data_out = 8'h37;
                    16'h63AD: data_out = 8'h36;
                    16'h63AE: data_out = 8'h35;
                    16'h63AF: data_out = 8'h34;
                    16'h63B0: data_out = 8'h33;
                    16'h63B1: data_out = 8'h32;
                    16'h63B2: data_out = 8'h31;
                    16'h63B3: data_out = 8'h30;
                    16'h63B4: data_out = 8'h2F;
                    16'h63B5: data_out = 8'h2E;
                    16'h63B6: data_out = 8'h2D;
                    16'h63B7: data_out = 8'h2C;
                    16'h63B8: data_out = 8'h2B;
                    16'h63B9: data_out = 8'h2A;
                    16'h63BA: data_out = 8'h29;
                    16'h63BB: data_out = 8'h28;
                    16'h63BC: data_out = 8'h27;
                    16'h63BD: data_out = 8'h26;
                    16'h63BE: data_out = 8'h25;
                    16'h63BF: data_out = 8'h24;
                    16'h63C0: data_out = 8'h23;
                    16'h63C1: data_out = 8'h22;
                    16'h63C2: data_out = 8'h21;
                    16'h63C3: data_out = 8'h20;
                    16'h63C4: data_out = 8'h1F;
                    16'h63C5: data_out = 8'h1E;
                    16'h63C6: data_out = 8'h1D;
                    16'h63C7: data_out = 8'h1C;
                    16'h63C8: data_out = 8'h1B;
                    16'h63C9: data_out = 8'h1A;
                    16'h63CA: data_out = 8'h19;
                    16'h63CB: data_out = 8'h18;
                    16'h63CC: data_out = 8'h17;
                    16'h63CD: data_out = 8'h16;
                    16'h63CE: data_out = 8'h15;
                    16'h63CF: data_out = 8'h14;
                    16'h63D0: data_out = 8'h13;
                    16'h63D1: data_out = 8'h12;
                    16'h63D2: data_out = 8'h11;
                    16'h63D3: data_out = 8'h10;
                    16'h63D4: data_out = 8'hF;
                    16'h63D5: data_out = 8'hE;
                    16'h63D6: data_out = 8'hD;
                    16'h63D7: data_out = 8'hC;
                    16'h63D8: data_out = 8'hB;
                    16'h63D9: data_out = 8'hA;
                    16'h63DA: data_out = 8'h9;
                    16'h63DB: data_out = 8'h8;
                    16'h63DC: data_out = 8'h7;
                    16'h63DD: data_out = 8'h6;
                    16'h63DE: data_out = 8'h5;
                    16'h63DF: data_out = 8'h4;
                    16'h63E0: data_out = 8'h3;
                    16'h63E1: data_out = 8'h2;
                    16'h63E2: data_out = 8'h1;
                    16'h63E3: data_out = 8'h0;
                    16'h63E4: data_out = 8'h81;
                    16'h63E5: data_out = 8'h82;
                    16'h63E6: data_out = 8'h83;
                    16'h63E7: data_out = 8'h84;
                    16'h63E8: data_out = 8'h85;
                    16'h63E9: data_out = 8'h86;
                    16'h63EA: data_out = 8'h87;
                    16'h63EB: data_out = 8'h88;
                    16'h63EC: data_out = 8'h89;
                    16'h63ED: data_out = 8'h8A;
                    16'h63EE: data_out = 8'h8B;
                    16'h63EF: data_out = 8'h8C;
                    16'h63F0: data_out = 8'h8D;
                    16'h63F1: data_out = 8'h8E;
                    16'h63F2: data_out = 8'h8F;
                    16'h63F3: data_out = 8'h90;
                    16'h63F4: data_out = 8'h91;
                    16'h63F5: data_out = 8'h92;
                    16'h63F6: data_out = 8'h93;
                    16'h63F7: data_out = 8'h94;
                    16'h63F8: data_out = 8'h95;
                    16'h63F9: data_out = 8'h96;
                    16'h63FA: data_out = 8'h97;
                    16'h63FB: data_out = 8'h98;
                    16'h63FC: data_out = 8'h99;
                    16'h63FD: data_out = 8'h9A;
                    16'h63FE: data_out = 8'h9B;
                    16'h63FF: data_out = 8'h9C;
                    16'h6400: data_out = 8'h64;
                    16'h6401: data_out = 8'h65;
                    16'h6402: data_out = 8'h66;
                    16'h6403: data_out = 8'h67;
                    16'h6404: data_out = 8'h68;
                    16'h6405: data_out = 8'h69;
                    16'h6406: data_out = 8'h6A;
                    16'h6407: data_out = 8'h6B;
                    16'h6408: data_out = 8'h6C;
                    16'h6409: data_out = 8'h6D;
                    16'h640A: data_out = 8'h6E;
                    16'h640B: data_out = 8'h6F;
                    16'h640C: data_out = 8'h70;
                    16'h640D: data_out = 8'h71;
                    16'h640E: data_out = 8'h72;
                    16'h640F: data_out = 8'h73;
                    16'h6410: data_out = 8'h74;
                    16'h6411: data_out = 8'h75;
                    16'h6412: data_out = 8'h76;
                    16'h6413: data_out = 8'h77;
                    16'h6414: data_out = 8'h78;
                    16'h6415: data_out = 8'h79;
                    16'h6416: data_out = 8'h7A;
                    16'h6417: data_out = 8'h7B;
                    16'h6418: data_out = 8'h7C;
                    16'h6419: data_out = 8'h7D;
                    16'h641A: data_out = 8'h7E;
                    16'h641B: data_out = 8'h7F;
                    16'h641C: data_out = 8'h80;
                    16'h641D: data_out = 8'h81;
                    16'h641E: data_out = 8'h82;
                    16'h641F: data_out = 8'h83;
                    16'h6420: data_out = 8'h84;
                    16'h6421: data_out = 8'h85;
                    16'h6422: data_out = 8'h86;
                    16'h6423: data_out = 8'h87;
                    16'h6424: data_out = 8'h88;
                    16'h6425: data_out = 8'h89;
                    16'h6426: data_out = 8'h8A;
                    16'h6427: data_out = 8'h8B;
                    16'h6428: data_out = 8'h8C;
                    16'h6429: data_out = 8'h8D;
                    16'h642A: data_out = 8'h8E;
                    16'h642B: data_out = 8'h8F;
                    16'h642C: data_out = 8'h90;
                    16'h642D: data_out = 8'h91;
                    16'h642E: data_out = 8'h92;
                    16'h642F: data_out = 8'h93;
                    16'h6430: data_out = 8'h94;
                    16'h6431: data_out = 8'h95;
                    16'h6432: data_out = 8'h96;
                    16'h6433: data_out = 8'h97;
                    16'h6434: data_out = 8'h98;
                    16'h6435: data_out = 8'h99;
                    16'h6436: data_out = 8'h9A;
                    16'h6437: data_out = 8'h9B;
                    16'h6438: data_out = 8'h9C;
                    16'h6439: data_out = 8'h9D;
                    16'h643A: data_out = 8'h9E;
                    16'h643B: data_out = 8'h9F;
                    16'h643C: data_out = 8'hA0;
                    16'h643D: data_out = 8'hA1;
                    16'h643E: data_out = 8'hA2;
                    16'h643F: data_out = 8'hA3;
                    16'h6440: data_out = 8'hA4;
                    16'h6441: data_out = 8'hA5;
                    16'h6442: data_out = 8'hA6;
                    16'h6443: data_out = 8'hA7;
                    16'h6444: data_out = 8'hA8;
                    16'h6445: data_out = 8'hA9;
                    16'h6446: data_out = 8'hAA;
                    16'h6447: data_out = 8'hAB;
                    16'h6448: data_out = 8'hAC;
                    16'h6449: data_out = 8'hAD;
                    16'h644A: data_out = 8'hAE;
                    16'h644B: data_out = 8'hAF;
                    16'h644C: data_out = 8'hB0;
                    16'h644D: data_out = 8'hB1;
                    16'h644E: data_out = 8'hB2;
                    16'h644F: data_out = 8'hB3;
                    16'h6450: data_out = 8'hB4;
                    16'h6451: data_out = 8'hB5;
                    16'h6452: data_out = 8'hB6;
                    16'h6453: data_out = 8'hB7;
                    16'h6454: data_out = 8'hB8;
                    16'h6455: data_out = 8'hB9;
                    16'h6456: data_out = 8'hBA;
                    16'h6457: data_out = 8'hBB;
                    16'h6458: data_out = 8'hBC;
                    16'h6459: data_out = 8'hBD;
                    16'h645A: data_out = 8'hBE;
                    16'h645B: data_out = 8'hBF;
                    16'h645C: data_out = 8'hC0;
                    16'h645D: data_out = 8'hC1;
                    16'h645E: data_out = 8'hC2;
                    16'h645F: data_out = 8'hC3;
                    16'h6460: data_out = 8'hC4;
                    16'h6461: data_out = 8'hC5;
                    16'h6462: data_out = 8'hC6;
                    16'h6463: data_out = 8'hC7;
                    16'h6464: data_out = 8'hC8;
                    16'h6465: data_out = 8'hC9;
                    16'h6466: data_out = 8'hCA;
                    16'h6467: data_out = 8'hCB;
                    16'h6468: data_out = 8'hCC;
                    16'h6469: data_out = 8'hCD;
                    16'h646A: data_out = 8'hCE;
                    16'h646B: data_out = 8'hCF;
                    16'h646C: data_out = 8'hD0;
                    16'h646D: data_out = 8'hD1;
                    16'h646E: data_out = 8'hD2;
                    16'h646F: data_out = 8'hD3;
                    16'h6470: data_out = 8'hD4;
                    16'h6471: data_out = 8'hD5;
                    16'h6472: data_out = 8'hD6;
                    16'h6473: data_out = 8'hD7;
                    16'h6474: data_out = 8'hD8;
                    16'h6475: data_out = 8'hD9;
                    16'h6476: data_out = 8'hDA;
                    16'h6477: data_out = 8'hDB;
                    16'h6478: data_out = 8'hDC;
                    16'h6479: data_out = 8'hDD;
                    16'h647A: data_out = 8'hDE;
                    16'h647B: data_out = 8'hDF;
                    16'h647C: data_out = 8'hE0;
                    16'h647D: data_out = 8'hE1;
                    16'h647E: data_out = 8'hE2;
                    16'h647F: data_out = 8'hE3;
                    16'h6480: data_out = 8'h64;
                    16'h6481: data_out = 8'h63;
                    16'h6482: data_out = 8'h62;
                    16'h6483: data_out = 8'h61;
                    16'h6484: data_out = 8'h60;
                    16'h6485: data_out = 8'h5F;
                    16'h6486: data_out = 8'h5E;
                    16'h6487: data_out = 8'h5D;
                    16'h6488: data_out = 8'h5C;
                    16'h6489: data_out = 8'h5B;
                    16'h648A: data_out = 8'h5A;
                    16'h648B: data_out = 8'h59;
                    16'h648C: data_out = 8'h58;
                    16'h648D: data_out = 8'h57;
                    16'h648E: data_out = 8'h56;
                    16'h648F: data_out = 8'h55;
                    16'h6490: data_out = 8'h54;
                    16'h6491: data_out = 8'h53;
                    16'h6492: data_out = 8'h52;
                    16'h6493: data_out = 8'h51;
                    16'h6494: data_out = 8'h50;
                    16'h6495: data_out = 8'h4F;
                    16'h6496: data_out = 8'h4E;
                    16'h6497: data_out = 8'h4D;
                    16'h6498: data_out = 8'h4C;
                    16'h6499: data_out = 8'h4B;
                    16'h649A: data_out = 8'h4A;
                    16'h649B: data_out = 8'h49;
                    16'h649C: data_out = 8'h48;
                    16'h649D: data_out = 8'h47;
                    16'h649E: data_out = 8'h46;
                    16'h649F: data_out = 8'h45;
                    16'h64A0: data_out = 8'h44;
                    16'h64A1: data_out = 8'h43;
                    16'h64A2: data_out = 8'h42;
                    16'h64A3: data_out = 8'h41;
                    16'h64A4: data_out = 8'h40;
                    16'h64A5: data_out = 8'h3F;
                    16'h64A6: data_out = 8'h3E;
                    16'h64A7: data_out = 8'h3D;
                    16'h64A8: data_out = 8'h3C;
                    16'h64A9: data_out = 8'h3B;
                    16'h64AA: data_out = 8'h3A;
                    16'h64AB: data_out = 8'h39;
                    16'h64AC: data_out = 8'h38;
                    16'h64AD: data_out = 8'h37;
                    16'h64AE: data_out = 8'h36;
                    16'h64AF: data_out = 8'h35;
                    16'h64B0: data_out = 8'h34;
                    16'h64B1: data_out = 8'h33;
                    16'h64B2: data_out = 8'h32;
                    16'h64B3: data_out = 8'h31;
                    16'h64B4: data_out = 8'h30;
                    16'h64B5: data_out = 8'h2F;
                    16'h64B6: data_out = 8'h2E;
                    16'h64B7: data_out = 8'h2D;
                    16'h64B8: data_out = 8'h2C;
                    16'h64B9: data_out = 8'h2B;
                    16'h64BA: data_out = 8'h2A;
                    16'h64BB: data_out = 8'h29;
                    16'h64BC: data_out = 8'h28;
                    16'h64BD: data_out = 8'h27;
                    16'h64BE: data_out = 8'h26;
                    16'h64BF: data_out = 8'h25;
                    16'h64C0: data_out = 8'h24;
                    16'h64C1: data_out = 8'h23;
                    16'h64C2: data_out = 8'h22;
                    16'h64C3: data_out = 8'h21;
                    16'h64C4: data_out = 8'h20;
                    16'h64C5: data_out = 8'h1F;
                    16'h64C6: data_out = 8'h1E;
                    16'h64C7: data_out = 8'h1D;
                    16'h64C8: data_out = 8'h1C;
                    16'h64C9: data_out = 8'h1B;
                    16'h64CA: data_out = 8'h1A;
                    16'h64CB: data_out = 8'h19;
                    16'h64CC: data_out = 8'h18;
                    16'h64CD: data_out = 8'h17;
                    16'h64CE: data_out = 8'h16;
                    16'h64CF: data_out = 8'h15;
                    16'h64D0: data_out = 8'h14;
                    16'h64D1: data_out = 8'h13;
                    16'h64D2: data_out = 8'h12;
                    16'h64D3: data_out = 8'h11;
                    16'h64D4: data_out = 8'h10;
                    16'h64D5: data_out = 8'hF;
                    16'h64D6: data_out = 8'hE;
                    16'h64D7: data_out = 8'hD;
                    16'h64D8: data_out = 8'hC;
                    16'h64D9: data_out = 8'hB;
                    16'h64DA: data_out = 8'hA;
                    16'h64DB: data_out = 8'h9;
                    16'h64DC: data_out = 8'h8;
                    16'h64DD: data_out = 8'h7;
                    16'h64DE: data_out = 8'h6;
                    16'h64DF: data_out = 8'h5;
                    16'h64E0: data_out = 8'h4;
                    16'h64E1: data_out = 8'h3;
                    16'h64E2: data_out = 8'h2;
                    16'h64E3: data_out = 8'h1;
                    16'h64E4: data_out = 8'h0;
                    16'h64E5: data_out = 8'h81;
                    16'h64E6: data_out = 8'h82;
                    16'h64E7: data_out = 8'h83;
                    16'h64E8: data_out = 8'h84;
                    16'h64E9: data_out = 8'h85;
                    16'h64EA: data_out = 8'h86;
                    16'h64EB: data_out = 8'h87;
                    16'h64EC: data_out = 8'h88;
                    16'h64ED: data_out = 8'h89;
                    16'h64EE: data_out = 8'h8A;
                    16'h64EF: data_out = 8'h8B;
                    16'h64F0: data_out = 8'h8C;
                    16'h64F1: data_out = 8'h8D;
                    16'h64F2: data_out = 8'h8E;
                    16'h64F3: data_out = 8'h8F;
                    16'h64F4: data_out = 8'h90;
                    16'h64F5: data_out = 8'h91;
                    16'h64F6: data_out = 8'h92;
                    16'h64F7: data_out = 8'h93;
                    16'h64F8: data_out = 8'h94;
                    16'h64F9: data_out = 8'h95;
                    16'h64FA: data_out = 8'h96;
                    16'h64FB: data_out = 8'h97;
                    16'h64FC: data_out = 8'h98;
                    16'h64FD: data_out = 8'h99;
                    16'h64FE: data_out = 8'h9A;
                    16'h64FF: data_out = 8'h9B;
                    16'h6500: data_out = 8'h65;
                    16'h6501: data_out = 8'h66;
                    16'h6502: data_out = 8'h67;
                    16'h6503: data_out = 8'h68;
                    16'h6504: data_out = 8'h69;
                    16'h6505: data_out = 8'h6A;
                    16'h6506: data_out = 8'h6B;
                    16'h6507: data_out = 8'h6C;
                    16'h6508: data_out = 8'h6D;
                    16'h6509: data_out = 8'h6E;
                    16'h650A: data_out = 8'h6F;
                    16'h650B: data_out = 8'h70;
                    16'h650C: data_out = 8'h71;
                    16'h650D: data_out = 8'h72;
                    16'h650E: data_out = 8'h73;
                    16'h650F: data_out = 8'h74;
                    16'h6510: data_out = 8'h75;
                    16'h6511: data_out = 8'h76;
                    16'h6512: data_out = 8'h77;
                    16'h6513: data_out = 8'h78;
                    16'h6514: data_out = 8'h79;
                    16'h6515: data_out = 8'h7A;
                    16'h6516: data_out = 8'h7B;
                    16'h6517: data_out = 8'h7C;
                    16'h6518: data_out = 8'h7D;
                    16'h6519: data_out = 8'h7E;
                    16'h651A: data_out = 8'h7F;
                    16'h651B: data_out = 8'h80;
                    16'h651C: data_out = 8'h81;
                    16'h651D: data_out = 8'h82;
                    16'h651E: data_out = 8'h83;
                    16'h651F: data_out = 8'h84;
                    16'h6520: data_out = 8'h85;
                    16'h6521: data_out = 8'h86;
                    16'h6522: data_out = 8'h87;
                    16'h6523: data_out = 8'h88;
                    16'h6524: data_out = 8'h89;
                    16'h6525: data_out = 8'h8A;
                    16'h6526: data_out = 8'h8B;
                    16'h6527: data_out = 8'h8C;
                    16'h6528: data_out = 8'h8D;
                    16'h6529: data_out = 8'h8E;
                    16'h652A: data_out = 8'h8F;
                    16'h652B: data_out = 8'h90;
                    16'h652C: data_out = 8'h91;
                    16'h652D: data_out = 8'h92;
                    16'h652E: data_out = 8'h93;
                    16'h652F: data_out = 8'h94;
                    16'h6530: data_out = 8'h95;
                    16'h6531: data_out = 8'h96;
                    16'h6532: data_out = 8'h97;
                    16'h6533: data_out = 8'h98;
                    16'h6534: data_out = 8'h99;
                    16'h6535: data_out = 8'h9A;
                    16'h6536: data_out = 8'h9B;
                    16'h6537: data_out = 8'h9C;
                    16'h6538: data_out = 8'h9D;
                    16'h6539: data_out = 8'h9E;
                    16'h653A: data_out = 8'h9F;
                    16'h653B: data_out = 8'hA0;
                    16'h653C: data_out = 8'hA1;
                    16'h653D: data_out = 8'hA2;
                    16'h653E: data_out = 8'hA3;
                    16'h653F: data_out = 8'hA4;
                    16'h6540: data_out = 8'hA5;
                    16'h6541: data_out = 8'hA6;
                    16'h6542: data_out = 8'hA7;
                    16'h6543: data_out = 8'hA8;
                    16'h6544: data_out = 8'hA9;
                    16'h6545: data_out = 8'hAA;
                    16'h6546: data_out = 8'hAB;
                    16'h6547: data_out = 8'hAC;
                    16'h6548: data_out = 8'hAD;
                    16'h6549: data_out = 8'hAE;
                    16'h654A: data_out = 8'hAF;
                    16'h654B: data_out = 8'hB0;
                    16'h654C: data_out = 8'hB1;
                    16'h654D: data_out = 8'hB2;
                    16'h654E: data_out = 8'hB3;
                    16'h654F: data_out = 8'hB4;
                    16'h6550: data_out = 8'hB5;
                    16'h6551: data_out = 8'hB6;
                    16'h6552: data_out = 8'hB7;
                    16'h6553: data_out = 8'hB8;
                    16'h6554: data_out = 8'hB9;
                    16'h6555: data_out = 8'hBA;
                    16'h6556: data_out = 8'hBB;
                    16'h6557: data_out = 8'hBC;
                    16'h6558: data_out = 8'hBD;
                    16'h6559: data_out = 8'hBE;
                    16'h655A: data_out = 8'hBF;
                    16'h655B: data_out = 8'hC0;
                    16'h655C: data_out = 8'hC1;
                    16'h655D: data_out = 8'hC2;
                    16'h655E: data_out = 8'hC3;
                    16'h655F: data_out = 8'hC4;
                    16'h6560: data_out = 8'hC5;
                    16'h6561: data_out = 8'hC6;
                    16'h6562: data_out = 8'hC7;
                    16'h6563: data_out = 8'hC8;
                    16'h6564: data_out = 8'hC9;
                    16'h6565: data_out = 8'hCA;
                    16'h6566: data_out = 8'hCB;
                    16'h6567: data_out = 8'hCC;
                    16'h6568: data_out = 8'hCD;
                    16'h6569: data_out = 8'hCE;
                    16'h656A: data_out = 8'hCF;
                    16'h656B: data_out = 8'hD0;
                    16'h656C: data_out = 8'hD1;
                    16'h656D: data_out = 8'hD2;
                    16'h656E: data_out = 8'hD3;
                    16'h656F: data_out = 8'hD4;
                    16'h6570: data_out = 8'hD5;
                    16'h6571: data_out = 8'hD6;
                    16'h6572: data_out = 8'hD7;
                    16'h6573: data_out = 8'hD8;
                    16'h6574: data_out = 8'hD9;
                    16'h6575: data_out = 8'hDA;
                    16'h6576: data_out = 8'hDB;
                    16'h6577: data_out = 8'hDC;
                    16'h6578: data_out = 8'hDD;
                    16'h6579: data_out = 8'hDE;
                    16'h657A: data_out = 8'hDF;
                    16'h657B: data_out = 8'hE0;
                    16'h657C: data_out = 8'hE1;
                    16'h657D: data_out = 8'hE2;
                    16'h657E: data_out = 8'hE3;
                    16'h657F: data_out = 8'hE4;
                    16'h6580: data_out = 8'h65;
                    16'h6581: data_out = 8'h64;
                    16'h6582: data_out = 8'h63;
                    16'h6583: data_out = 8'h62;
                    16'h6584: data_out = 8'h61;
                    16'h6585: data_out = 8'h60;
                    16'h6586: data_out = 8'h5F;
                    16'h6587: data_out = 8'h5E;
                    16'h6588: data_out = 8'h5D;
                    16'h6589: data_out = 8'h5C;
                    16'h658A: data_out = 8'h5B;
                    16'h658B: data_out = 8'h5A;
                    16'h658C: data_out = 8'h59;
                    16'h658D: data_out = 8'h58;
                    16'h658E: data_out = 8'h57;
                    16'h658F: data_out = 8'h56;
                    16'h6590: data_out = 8'h55;
                    16'h6591: data_out = 8'h54;
                    16'h6592: data_out = 8'h53;
                    16'h6593: data_out = 8'h52;
                    16'h6594: data_out = 8'h51;
                    16'h6595: data_out = 8'h50;
                    16'h6596: data_out = 8'h4F;
                    16'h6597: data_out = 8'h4E;
                    16'h6598: data_out = 8'h4D;
                    16'h6599: data_out = 8'h4C;
                    16'h659A: data_out = 8'h4B;
                    16'h659B: data_out = 8'h4A;
                    16'h659C: data_out = 8'h49;
                    16'h659D: data_out = 8'h48;
                    16'h659E: data_out = 8'h47;
                    16'h659F: data_out = 8'h46;
                    16'h65A0: data_out = 8'h45;
                    16'h65A1: data_out = 8'h44;
                    16'h65A2: data_out = 8'h43;
                    16'h65A3: data_out = 8'h42;
                    16'h65A4: data_out = 8'h41;
                    16'h65A5: data_out = 8'h40;
                    16'h65A6: data_out = 8'h3F;
                    16'h65A7: data_out = 8'h3E;
                    16'h65A8: data_out = 8'h3D;
                    16'h65A9: data_out = 8'h3C;
                    16'h65AA: data_out = 8'h3B;
                    16'h65AB: data_out = 8'h3A;
                    16'h65AC: data_out = 8'h39;
                    16'h65AD: data_out = 8'h38;
                    16'h65AE: data_out = 8'h37;
                    16'h65AF: data_out = 8'h36;
                    16'h65B0: data_out = 8'h35;
                    16'h65B1: data_out = 8'h34;
                    16'h65B2: data_out = 8'h33;
                    16'h65B3: data_out = 8'h32;
                    16'h65B4: data_out = 8'h31;
                    16'h65B5: data_out = 8'h30;
                    16'h65B6: data_out = 8'h2F;
                    16'h65B7: data_out = 8'h2E;
                    16'h65B8: data_out = 8'h2D;
                    16'h65B9: data_out = 8'h2C;
                    16'h65BA: data_out = 8'h2B;
                    16'h65BB: data_out = 8'h2A;
                    16'h65BC: data_out = 8'h29;
                    16'h65BD: data_out = 8'h28;
                    16'h65BE: data_out = 8'h27;
                    16'h65BF: data_out = 8'h26;
                    16'h65C0: data_out = 8'h25;
                    16'h65C1: data_out = 8'h24;
                    16'h65C2: data_out = 8'h23;
                    16'h65C3: data_out = 8'h22;
                    16'h65C4: data_out = 8'h21;
                    16'h65C5: data_out = 8'h20;
                    16'h65C6: data_out = 8'h1F;
                    16'h65C7: data_out = 8'h1E;
                    16'h65C8: data_out = 8'h1D;
                    16'h65C9: data_out = 8'h1C;
                    16'h65CA: data_out = 8'h1B;
                    16'h65CB: data_out = 8'h1A;
                    16'h65CC: data_out = 8'h19;
                    16'h65CD: data_out = 8'h18;
                    16'h65CE: data_out = 8'h17;
                    16'h65CF: data_out = 8'h16;
                    16'h65D0: data_out = 8'h15;
                    16'h65D1: data_out = 8'h14;
                    16'h65D2: data_out = 8'h13;
                    16'h65D3: data_out = 8'h12;
                    16'h65D4: data_out = 8'h11;
                    16'h65D5: data_out = 8'h10;
                    16'h65D6: data_out = 8'hF;
                    16'h65D7: data_out = 8'hE;
                    16'h65D8: data_out = 8'hD;
                    16'h65D9: data_out = 8'hC;
                    16'h65DA: data_out = 8'hB;
                    16'h65DB: data_out = 8'hA;
                    16'h65DC: data_out = 8'h9;
                    16'h65DD: data_out = 8'h8;
                    16'h65DE: data_out = 8'h7;
                    16'h65DF: data_out = 8'h6;
                    16'h65E0: data_out = 8'h5;
                    16'h65E1: data_out = 8'h4;
                    16'h65E2: data_out = 8'h3;
                    16'h65E3: data_out = 8'h2;
                    16'h65E4: data_out = 8'h1;
                    16'h65E5: data_out = 8'h0;
                    16'h65E6: data_out = 8'h81;
                    16'h65E7: data_out = 8'h82;
                    16'h65E8: data_out = 8'h83;
                    16'h65E9: data_out = 8'h84;
                    16'h65EA: data_out = 8'h85;
                    16'h65EB: data_out = 8'h86;
                    16'h65EC: data_out = 8'h87;
                    16'h65ED: data_out = 8'h88;
                    16'h65EE: data_out = 8'h89;
                    16'h65EF: data_out = 8'h8A;
                    16'h65F0: data_out = 8'h8B;
                    16'h65F1: data_out = 8'h8C;
                    16'h65F2: data_out = 8'h8D;
                    16'h65F3: data_out = 8'h8E;
                    16'h65F4: data_out = 8'h8F;
                    16'h65F5: data_out = 8'h90;
                    16'h65F6: data_out = 8'h91;
                    16'h65F7: data_out = 8'h92;
                    16'h65F8: data_out = 8'h93;
                    16'h65F9: data_out = 8'h94;
                    16'h65FA: data_out = 8'h95;
                    16'h65FB: data_out = 8'h96;
                    16'h65FC: data_out = 8'h97;
                    16'h65FD: data_out = 8'h98;
                    16'h65FE: data_out = 8'h99;
                    16'h65FF: data_out = 8'h9A;
                    16'h6600: data_out = 8'h66;
                    16'h6601: data_out = 8'h67;
                    16'h6602: data_out = 8'h68;
                    16'h6603: data_out = 8'h69;
                    16'h6604: data_out = 8'h6A;
                    16'h6605: data_out = 8'h6B;
                    16'h6606: data_out = 8'h6C;
                    16'h6607: data_out = 8'h6D;
                    16'h6608: data_out = 8'h6E;
                    16'h6609: data_out = 8'h6F;
                    16'h660A: data_out = 8'h70;
                    16'h660B: data_out = 8'h71;
                    16'h660C: data_out = 8'h72;
                    16'h660D: data_out = 8'h73;
                    16'h660E: data_out = 8'h74;
                    16'h660F: data_out = 8'h75;
                    16'h6610: data_out = 8'h76;
                    16'h6611: data_out = 8'h77;
                    16'h6612: data_out = 8'h78;
                    16'h6613: data_out = 8'h79;
                    16'h6614: data_out = 8'h7A;
                    16'h6615: data_out = 8'h7B;
                    16'h6616: data_out = 8'h7C;
                    16'h6617: data_out = 8'h7D;
                    16'h6618: data_out = 8'h7E;
                    16'h6619: data_out = 8'h7F;
                    16'h661A: data_out = 8'h80;
                    16'h661B: data_out = 8'h81;
                    16'h661C: data_out = 8'h82;
                    16'h661D: data_out = 8'h83;
                    16'h661E: data_out = 8'h84;
                    16'h661F: data_out = 8'h85;
                    16'h6620: data_out = 8'h86;
                    16'h6621: data_out = 8'h87;
                    16'h6622: data_out = 8'h88;
                    16'h6623: data_out = 8'h89;
                    16'h6624: data_out = 8'h8A;
                    16'h6625: data_out = 8'h8B;
                    16'h6626: data_out = 8'h8C;
                    16'h6627: data_out = 8'h8D;
                    16'h6628: data_out = 8'h8E;
                    16'h6629: data_out = 8'h8F;
                    16'h662A: data_out = 8'h90;
                    16'h662B: data_out = 8'h91;
                    16'h662C: data_out = 8'h92;
                    16'h662D: data_out = 8'h93;
                    16'h662E: data_out = 8'h94;
                    16'h662F: data_out = 8'h95;
                    16'h6630: data_out = 8'h96;
                    16'h6631: data_out = 8'h97;
                    16'h6632: data_out = 8'h98;
                    16'h6633: data_out = 8'h99;
                    16'h6634: data_out = 8'h9A;
                    16'h6635: data_out = 8'h9B;
                    16'h6636: data_out = 8'h9C;
                    16'h6637: data_out = 8'h9D;
                    16'h6638: data_out = 8'h9E;
                    16'h6639: data_out = 8'h9F;
                    16'h663A: data_out = 8'hA0;
                    16'h663B: data_out = 8'hA1;
                    16'h663C: data_out = 8'hA2;
                    16'h663D: data_out = 8'hA3;
                    16'h663E: data_out = 8'hA4;
                    16'h663F: data_out = 8'hA5;
                    16'h6640: data_out = 8'hA6;
                    16'h6641: data_out = 8'hA7;
                    16'h6642: data_out = 8'hA8;
                    16'h6643: data_out = 8'hA9;
                    16'h6644: data_out = 8'hAA;
                    16'h6645: data_out = 8'hAB;
                    16'h6646: data_out = 8'hAC;
                    16'h6647: data_out = 8'hAD;
                    16'h6648: data_out = 8'hAE;
                    16'h6649: data_out = 8'hAF;
                    16'h664A: data_out = 8'hB0;
                    16'h664B: data_out = 8'hB1;
                    16'h664C: data_out = 8'hB2;
                    16'h664D: data_out = 8'hB3;
                    16'h664E: data_out = 8'hB4;
                    16'h664F: data_out = 8'hB5;
                    16'h6650: data_out = 8'hB6;
                    16'h6651: data_out = 8'hB7;
                    16'h6652: data_out = 8'hB8;
                    16'h6653: data_out = 8'hB9;
                    16'h6654: data_out = 8'hBA;
                    16'h6655: data_out = 8'hBB;
                    16'h6656: data_out = 8'hBC;
                    16'h6657: data_out = 8'hBD;
                    16'h6658: data_out = 8'hBE;
                    16'h6659: data_out = 8'hBF;
                    16'h665A: data_out = 8'hC0;
                    16'h665B: data_out = 8'hC1;
                    16'h665C: data_out = 8'hC2;
                    16'h665D: data_out = 8'hC3;
                    16'h665E: data_out = 8'hC4;
                    16'h665F: data_out = 8'hC5;
                    16'h6660: data_out = 8'hC6;
                    16'h6661: data_out = 8'hC7;
                    16'h6662: data_out = 8'hC8;
                    16'h6663: data_out = 8'hC9;
                    16'h6664: data_out = 8'hCA;
                    16'h6665: data_out = 8'hCB;
                    16'h6666: data_out = 8'hCC;
                    16'h6667: data_out = 8'hCD;
                    16'h6668: data_out = 8'hCE;
                    16'h6669: data_out = 8'hCF;
                    16'h666A: data_out = 8'hD0;
                    16'h666B: data_out = 8'hD1;
                    16'h666C: data_out = 8'hD2;
                    16'h666D: data_out = 8'hD3;
                    16'h666E: data_out = 8'hD4;
                    16'h666F: data_out = 8'hD5;
                    16'h6670: data_out = 8'hD6;
                    16'h6671: data_out = 8'hD7;
                    16'h6672: data_out = 8'hD8;
                    16'h6673: data_out = 8'hD9;
                    16'h6674: data_out = 8'hDA;
                    16'h6675: data_out = 8'hDB;
                    16'h6676: data_out = 8'hDC;
                    16'h6677: data_out = 8'hDD;
                    16'h6678: data_out = 8'hDE;
                    16'h6679: data_out = 8'hDF;
                    16'h667A: data_out = 8'hE0;
                    16'h667B: data_out = 8'hE1;
                    16'h667C: data_out = 8'hE2;
                    16'h667D: data_out = 8'hE3;
                    16'h667E: data_out = 8'hE4;
                    16'h667F: data_out = 8'hE5;
                    16'h6680: data_out = 8'h66;
                    16'h6681: data_out = 8'h65;
                    16'h6682: data_out = 8'h64;
                    16'h6683: data_out = 8'h63;
                    16'h6684: data_out = 8'h62;
                    16'h6685: data_out = 8'h61;
                    16'h6686: data_out = 8'h60;
                    16'h6687: data_out = 8'h5F;
                    16'h6688: data_out = 8'h5E;
                    16'h6689: data_out = 8'h5D;
                    16'h668A: data_out = 8'h5C;
                    16'h668B: data_out = 8'h5B;
                    16'h668C: data_out = 8'h5A;
                    16'h668D: data_out = 8'h59;
                    16'h668E: data_out = 8'h58;
                    16'h668F: data_out = 8'h57;
                    16'h6690: data_out = 8'h56;
                    16'h6691: data_out = 8'h55;
                    16'h6692: data_out = 8'h54;
                    16'h6693: data_out = 8'h53;
                    16'h6694: data_out = 8'h52;
                    16'h6695: data_out = 8'h51;
                    16'h6696: data_out = 8'h50;
                    16'h6697: data_out = 8'h4F;
                    16'h6698: data_out = 8'h4E;
                    16'h6699: data_out = 8'h4D;
                    16'h669A: data_out = 8'h4C;
                    16'h669B: data_out = 8'h4B;
                    16'h669C: data_out = 8'h4A;
                    16'h669D: data_out = 8'h49;
                    16'h669E: data_out = 8'h48;
                    16'h669F: data_out = 8'h47;
                    16'h66A0: data_out = 8'h46;
                    16'h66A1: data_out = 8'h45;
                    16'h66A2: data_out = 8'h44;
                    16'h66A3: data_out = 8'h43;
                    16'h66A4: data_out = 8'h42;
                    16'h66A5: data_out = 8'h41;
                    16'h66A6: data_out = 8'h40;
                    16'h66A7: data_out = 8'h3F;
                    16'h66A8: data_out = 8'h3E;
                    16'h66A9: data_out = 8'h3D;
                    16'h66AA: data_out = 8'h3C;
                    16'h66AB: data_out = 8'h3B;
                    16'h66AC: data_out = 8'h3A;
                    16'h66AD: data_out = 8'h39;
                    16'h66AE: data_out = 8'h38;
                    16'h66AF: data_out = 8'h37;
                    16'h66B0: data_out = 8'h36;
                    16'h66B1: data_out = 8'h35;
                    16'h66B2: data_out = 8'h34;
                    16'h66B3: data_out = 8'h33;
                    16'h66B4: data_out = 8'h32;
                    16'h66B5: data_out = 8'h31;
                    16'h66B6: data_out = 8'h30;
                    16'h66B7: data_out = 8'h2F;
                    16'h66B8: data_out = 8'h2E;
                    16'h66B9: data_out = 8'h2D;
                    16'h66BA: data_out = 8'h2C;
                    16'h66BB: data_out = 8'h2B;
                    16'h66BC: data_out = 8'h2A;
                    16'h66BD: data_out = 8'h29;
                    16'h66BE: data_out = 8'h28;
                    16'h66BF: data_out = 8'h27;
                    16'h66C0: data_out = 8'h26;
                    16'h66C1: data_out = 8'h25;
                    16'h66C2: data_out = 8'h24;
                    16'h66C3: data_out = 8'h23;
                    16'h66C4: data_out = 8'h22;
                    16'h66C5: data_out = 8'h21;
                    16'h66C6: data_out = 8'h20;
                    16'h66C7: data_out = 8'h1F;
                    16'h66C8: data_out = 8'h1E;
                    16'h66C9: data_out = 8'h1D;
                    16'h66CA: data_out = 8'h1C;
                    16'h66CB: data_out = 8'h1B;
                    16'h66CC: data_out = 8'h1A;
                    16'h66CD: data_out = 8'h19;
                    16'h66CE: data_out = 8'h18;
                    16'h66CF: data_out = 8'h17;
                    16'h66D0: data_out = 8'h16;
                    16'h66D1: data_out = 8'h15;
                    16'h66D2: data_out = 8'h14;
                    16'h66D3: data_out = 8'h13;
                    16'h66D4: data_out = 8'h12;
                    16'h66D5: data_out = 8'h11;
                    16'h66D6: data_out = 8'h10;
                    16'h66D7: data_out = 8'hF;
                    16'h66D8: data_out = 8'hE;
                    16'h66D9: data_out = 8'hD;
                    16'h66DA: data_out = 8'hC;
                    16'h66DB: data_out = 8'hB;
                    16'h66DC: data_out = 8'hA;
                    16'h66DD: data_out = 8'h9;
                    16'h66DE: data_out = 8'h8;
                    16'h66DF: data_out = 8'h7;
                    16'h66E0: data_out = 8'h6;
                    16'h66E1: data_out = 8'h5;
                    16'h66E2: data_out = 8'h4;
                    16'h66E3: data_out = 8'h3;
                    16'h66E4: data_out = 8'h2;
                    16'h66E5: data_out = 8'h1;
                    16'h66E6: data_out = 8'h0;
                    16'h66E7: data_out = 8'h81;
                    16'h66E8: data_out = 8'h82;
                    16'h66E9: data_out = 8'h83;
                    16'h66EA: data_out = 8'h84;
                    16'h66EB: data_out = 8'h85;
                    16'h66EC: data_out = 8'h86;
                    16'h66ED: data_out = 8'h87;
                    16'h66EE: data_out = 8'h88;
                    16'h66EF: data_out = 8'h89;
                    16'h66F0: data_out = 8'h8A;
                    16'h66F1: data_out = 8'h8B;
                    16'h66F2: data_out = 8'h8C;
                    16'h66F3: data_out = 8'h8D;
                    16'h66F4: data_out = 8'h8E;
                    16'h66F5: data_out = 8'h8F;
                    16'h66F6: data_out = 8'h90;
                    16'h66F7: data_out = 8'h91;
                    16'h66F8: data_out = 8'h92;
                    16'h66F9: data_out = 8'h93;
                    16'h66FA: data_out = 8'h94;
                    16'h66FB: data_out = 8'h95;
                    16'h66FC: data_out = 8'h96;
                    16'h66FD: data_out = 8'h97;
                    16'h66FE: data_out = 8'h98;
                    16'h66FF: data_out = 8'h99;
                    16'h6700: data_out = 8'h67;
                    16'h6701: data_out = 8'h68;
                    16'h6702: data_out = 8'h69;
                    16'h6703: data_out = 8'h6A;
                    16'h6704: data_out = 8'h6B;
                    16'h6705: data_out = 8'h6C;
                    16'h6706: data_out = 8'h6D;
                    16'h6707: data_out = 8'h6E;
                    16'h6708: data_out = 8'h6F;
                    16'h6709: data_out = 8'h70;
                    16'h670A: data_out = 8'h71;
                    16'h670B: data_out = 8'h72;
                    16'h670C: data_out = 8'h73;
                    16'h670D: data_out = 8'h74;
                    16'h670E: data_out = 8'h75;
                    16'h670F: data_out = 8'h76;
                    16'h6710: data_out = 8'h77;
                    16'h6711: data_out = 8'h78;
                    16'h6712: data_out = 8'h79;
                    16'h6713: data_out = 8'h7A;
                    16'h6714: data_out = 8'h7B;
                    16'h6715: data_out = 8'h7C;
                    16'h6716: data_out = 8'h7D;
                    16'h6717: data_out = 8'h7E;
                    16'h6718: data_out = 8'h7F;
                    16'h6719: data_out = 8'h80;
                    16'h671A: data_out = 8'h81;
                    16'h671B: data_out = 8'h82;
                    16'h671C: data_out = 8'h83;
                    16'h671D: data_out = 8'h84;
                    16'h671E: data_out = 8'h85;
                    16'h671F: data_out = 8'h86;
                    16'h6720: data_out = 8'h87;
                    16'h6721: data_out = 8'h88;
                    16'h6722: data_out = 8'h89;
                    16'h6723: data_out = 8'h8A;
                    16'h6724: data_out = 8'h8B;
                    16'h6725: data_out = 8'h8C;
                    16'h6726: data_out = 8'h8D;
                    16'h6727: data_out = 8'h8E;
                    16'h6728: data_out = 8'h8F;
                    16'h6729: data_out = 8'h90;
                    16'h672A: data_out = 8'h91;
                    16'h672B: data_out = 8'h92;
                    16'h672C: data_out = 8'h93;
                    16'h672D: data_out = 8'h94;
                    16'h672E: data_out = 8'h95;
                    16'h672F: data_out = 8'h96;
                    16'h6730: data_out = 8'h97;
                    16'h6731: data_out = 8'h98;
                    16'h6732: data_out = 8'h99;
                    16'h6733: data_out = 8'h9A;
                    16'h6734: data_out = 8'h9B;
                    16'h6735: data_out = 8'h9C;
                    16'h6736: data_out = 8'h9D;
                    16'h6737: data_out = 8'h9E;
                    16'h6738: data_out = 8'h9F;
                    16'h6739: data_out = 8'hA0;
                    16'h673A: data_out = 8'hA1;
                    16'h673B: data_out = 8'hA2;
                    16'h673C: data_out = 8'hA3;
                    16'h673D: data_out = 8'hA4;
                    16'h673E: data_out = 8'hA5;
                    16'h673F: data_out = 8'hA6;
                    16'h6740: data_out = 8'hA7;
                    16'h6741: data_out = 8'hA8;
                    16'h6742: data_out = 8'hA9;
                    16'h6743: data_out = 8'hAA;
                    16'h6744: data_out = 8'hAB;
                    16'h6745: data_out = 8'hAC;
                    16'h6746: data_out = 8'hAD;
                    16'h6747: data_out = 8'hAE;
                    16'h6748: data_out = 8'hAF;
                    16'h6749: data_out = 8'hB0;
                    16'h674A: data_out = 8'hB1;
                    16'h674B: data_out = 8'hB2;
                    16'h674C: data_out = 8'hB3;
                    16'h674D: data_out = 8'hB4;
                    16'h674E: data_out = 8'hB5;
                    16'h674F: data_out = 8'hB6;
                    16'h6750: data_out = 8'hB7;
                    16'h6751: data_out = 8'hB8;
                    16'h6752: data_out = 8'hB9;
                    16'h6753: data_out = 8'hBA;
                    16'h6754: data_out = 8'hBB;
                    16'h6755: data_out = 8'hBC;
                    16'h6756: data_out = 8'hBD;
                    16'h6757: data_out = 8'hBE;
                    16'h6758: data_out = 8'hBF;
                    16'h6759: data_out = 8'hC0;
                    16'h675A: data_out = 8'hC1;
                    16'h675B: data_out = 8'hC2;
                    16'h675C: data_out = 8'hC3;
                    16'h675D: data_out = 8'hC4;
                    16'h675E: data_out = 8'hC5;
                    16'h675F: data_out = 8'hC6;
                    16'h6760: data_out = 8'hC7;
                    16'h6761: data_out = 8'hC8;
                    16'h6762: data_out = 8'hC9;
                    16'h6763: data_out = 8'hCA;
                    16'h6764: data_out = 8'hCB;
                    16'h6765: data_out = 8'hCC;
                    16'h6766: data_out = 8'hCD;
                    16'h6767: data_out = 8'hCE;
                    16'h6768: data_out = 8'hCF;
                    16'h6769: data_out = 8'hD0;
                    16'h676A: data_out = 8'hD1;
                    16'h676B: data_out = 8'hD2;
                    16'h676C: data_out = 8'hD3;
                    16'h676D: data_out = 8'hD4;
                    16'h676E: data_out = 8'hD5;
                    16'h676F: data_out = 8'hD6;
                    16'h6770: data_out = 8'hD7;
                    16'h6771: data_out = 8'hD8;
                    16'h6772: data_out = 8'hD9;
                    16'h6773: data_out = 8'hDA;
                    16'h6774: data_out = 8'hDB;
                    16'h6775: data_out = 8'hDC;
                    16'h6776: data_out = 8'hDD;
                    16'h6777: data_out = 8'hDE;
                    16'h6778: data_out = 8'hDF;
                    16'h6779: data_out = 8'hE0;
                    16'h677A: data_out = 8'hE1;
                    16'h677B: data_out = 8'hE2;
                    16'h677C: data_out = 8'hE3;
                    16'h677D: data_out = 8'hE4;
                    16'h677E: data_out = 8'hE5;
                    16'h677F: data_out = 8'hE6;
                    16'h6780: data_out = 8'h67;
                    16'h6781: data_out = 8'h66;
                    16'h6782: data_out = 8'h65;
                    16'h6783: data_out = 8'h64;
                    16'h6784: data_out = 8'h63;
                    16'h6785: data_out = 8'h62;
                    16'h6786: data_out = 8'h61;
                    16'h6787: data_out = 8'h60;
                    16'h6788: data_out = 8'h5F;
                    16'h6789: data_out = 8'h5E;
                    16'h678A: data_out = 8'h5D;
                    16'h678B: data_out = 8'h5C;
                    16'h678C: data_out = 8'h5B;
                    16'h678D: data_out = 8'h5A;
                    16'h678E: data_out = 8'h59;
                    16'h678F: data_out = 8'h58;
                    16'h6790: data_out = 8'h57;
                    16'h6791: data_out = 8'h56;
                    16'h6792: data_out = 8'h55;
                    16'h6793: data_out = 8'h54;
                    16'h6794: data_out = 8'h53;
                    16'h6795: data_out = 8'h52;
                    16'h6796: data_out = 8'h51;
                    16'h6797: data_out = 8'h50;
                    16'h6798: data_out = 8'h4F;
                    16'h6799: data_out = 8'h4E;
                    16'h679A: data_out = 8'h4D;
                    16'h679B: data_out = 8'h4C;
                    16'h679C: data_out = 8'h4B;
                    16'h679D: data_out = 8'h4A;
                    16'h679E: data_out = 8'h49;
                    16'h679F: data_out = 8'h48;
                    16'h67A0: data_out = 8'h47;
                    16'h67A1: data_out = 8'h46;
                    16'h67A2: data_out = 8'h45;
                    16'h67A3: data_out = 8'h44;
                    16'h67A4: data_out = 8'h43;
                    16'h67A5: data_out = 8'h42;
                    16'h67A6: data_out = 8'h41;
                    16'h67A7: data_out = 8'h40;
                    16'h67A8: data_out = 8'h3F;
                    16'h67A9: data_out = 8'h3E;
                    16'h67AA: data_out = 8'h3D;
                    16'h67AB: data_out = 8'h3C;
                    16'h67AC: data_out = 8'h3B;
                    16'h67AD: data_out = 8'h3A;
                    16'h67AE: data_out = 8'h39;
                    16'h67AF: data_out = 8'h38;
                    16'h67B0: data_out = 8'h37;
                    16'h67B1: data_out = 8'h36;
                    16'h67B2: data_out = 8'h35;
                    16'h67B3: data_out = 8'h34;
                    16'h67B4: data_out = 8'h33;
                    16'h67B5: data_out = 8'h32;
                    16'h67B6: data_out = 8'h31;
                    16'h67B7: data_out = 8'h30;
                    16'h67B8: data_out = 8'h2F;
                    16'h67B9: data_out = 8'h2E;
                    16'h67BA: data_out = 8'h2D;
                    16'h67BB: data_out = 8'h2C;
                    16'h67BC: data_out = 8'h2B;
                    16'h67BD: data_out = 8'h2A;
                    16'h67BE: data_out = 8'h29;
                    16'h67BF: data_out = 8'h28;
                    16'h67C0: data_out = 8'h27;
                    16'h67C1: data_out = 8'h26;
                    16'h67C2: data_out = 8'h25;
                    16'h67C3: data_out = 8'h24;
                    16'h67C4: data_out = 8'h23;
                    16'h67C5: data_out = 8'h22;
                    16'h67C6: data_out = 8'h21;
                    16'h67C7: data_out = 8'h20;
                    16'h67C8: data_out = 8'h1F;
                    16'h67C9: data_out = 8'h1E;
                    16'h67CA: data_out = 8'h1D;
                    16'h67CB: data_out = 8'h1C;
                    16'h67CC: data_out = 8'h1B;
                    16'h67CD: data_out = 8'h1A;
                    16'h67CE: data_out = 8'h19;
                    16'h67CF: data_out = 8'h18;
                    16'h67D0: data_out = 8'h17;
                    16'h67D1: data_out = 8'h16;
                    16'h67D2: data_out = 8'h15;
                    16'h67D3: data_out = 8'h14;
                    16'h67D4: data_out = 8'h13;
                    16'h67D5: data_out = 8'h12;
                    16'h67D6: data_out = 8'h11;
                    16'h67D7: data_out = 8'h10;
                    16'h67D8: data_out = 8'hF;
                    16'h67D9: data_out = 8'hE;
                    16'h67DA: data_out = 8'hD;
                    16'h67DB: data_out = 8'hC;
                    16'h67DC: data_out = 8'hB;
                    16'h67DD: data_out = 8'hA;
                    16'h67DE: data_out = 8'h9;
                    16'h67DF: data_out = 8'h8;
                    16'h67E0: data_out = 8'h7;
                    16'h67E1: data_out = 8'h6;
                    16'h67E2: data_out = 8'h5;
                    16'h67E3: data_out = 8'h4;
                    16'h67E4: data_out = 8'h3;
                    16'h67E5: data_out = 8'h2;
                    16'h67E6: data_out = 8'h1;
                    16'h67E7: data_out = 8'h0;
                    16'h67E8: data_out = 8'h81;
                    16'h67E9: data_out = 8'h82;
                    16'h67EA: data_out = 8'h83;
                    16'h67EB: data_out = 8'h84;
                    16'h67EC: data_out = 8'h85;
                    16'h67ED: data_out = 8'h86;
                    16'h67EE: data_out = 8'h87;
                    16'h67EF: data_out = 8'h88;
                    16'h67F0: data_out = 8'h89;
                    16'h67F1: data_out = 8'h8A;
                    16'h67F2: data_out = 8'h8B;
                    16'h67F3: data_out = 8'h8C;
                    16'h67F4: data_out = 8'h8D;
                    16'h67F5: data_out = 8'h8E;
                    16'h67F6: data_out = 8'h8F;
                    16'h67F7: data_out = 8'h90;
                    16'h67F8: data_out = 8'h91;
                    16'h67F9: data_out = 8'h92;
                    16'h67FA: data_out = 8'h93;
                    16'h67FB: data_out = 8'h94;
                    16'h67FC: data_out = 8'h95;
                    16'h67FD: data_out = 8'h96;
                    16'h67FE: data_out = 8'h97;
                    16'h67FF: data_out = 8'h98;
                    16'h6800: data_out = 8'h68;
                    16'h6801: data_out = 8'h69;
                    16'h6802: data_out = 8'h6A;
                    16'h6803: data_out = 8'h6B;
                    16'h6804: data_out = 8'h6C;
                    16'h6805: data_out = 8'h6D;
                    16'h6806: data_out = 8'h6E;
                    16'h6807: data_out = 8'h6F;
                    16'h6808: data_out = 8'h70;
                    16'h6809: data_out = 8'h71;
                    16'h680A: data_out = 8'h72;
                    16'h680B: data_out = 8'h73;
                    16'h680C: data_out = 8'h74;
                    16'h680D: data_out = 8'h75;
                    16'h680E: data_out = 8'h76;
                    16'h680F: data_out = 8'h77;
                    16'h6810: data_out = 8'h78;
                    16'h6811: data_out = 8'h79;
                    16'h6812: data_out = 8'h7A;
                    16'h6813: data_out = 8'h7B;
                    16'h6814: data_out = 8'h7C;
                    16'h6815: data_out = 8'h7D;
                    16'h6816: data_out = 8'h7E;
                    16'h6817: data_out = 8'h7F;
                    16'h6818: data_out = 8'h80;
                    16'h6819: data_out = 8'h81;
                    16'h681A: data_out = 8'h82;
                    16'h681B: data_out = 8'h83;
                    16'h681C: data_out = 8'h84;
                    16'h681D: data_out = 8'h85;
                    16'h681E: data_out = 8'h86;
                    16'h681F: data_out = 8'h87;
                    16'h6820: data_out = 8'h88;
                    16'h6821: data_out = 8'h89;
                    16'h6822: data_out = 8'h8A;
                    16'h6823: data_out = 8'h8B;
                    16'h6824: data_out = 8'h8C;
                    16'h6825: data_out = 8'h8D;
                    16'h6826: data_out = 8'h8E;
                    16'h6827: data_out = 8'h8F;
                    16'h6828: data_out = 8'h90;
                    16'h6829: data_out = 8'h91;
                    16'h682A: data_out = 8'h92;
                    16'h682B: data_out = 8'h93;
                    16'h682C: data_out = 8'h94;
                    16'h682D: data_out = 8'h95;
                    16'h682E: data_out = 8'h96;
                    16'h682F: data_out = 8'h97;
                    16'h6830: data_out = 8'h98;
                    16'h6831: data_out = 8'h99;
                    16'h6832: data_out = 8'h9A;
                    16'h6833: data_out = 8'h9B;
                    16'h6834: data_out = 8'h9C;
                    16'h6835: data_out = 8'h9D;
                    16'h6836: data_out = 8'h9E;
                    16'h6837: data_out = 8'h9F;
                    16'h6838: data_out = 8'hA0;
                    16'h6839: data_out = 8'hA1;
                    16'h683A: data_out = 8'hA2;
                    16'h683B: data_out = 8'hA3;
                    16'h683C: data_out = 8'hA4;
                    16'h683D: data_out = 8'hA5;
                    16'h683E: data_out = 8'hA6;
                    16'h683F: data_out = 8'hA7;
                    16'h6840: data_out = 8'hA8;
                    16'h6841: data_out = 8'hA9;
                    16'h6842: data_out = 8'hAA;
                    16'h6843: data_out = 8'hAB;
                    16'h6844: data_out = 8'hAC;
                    16'h6845: data_out = 8'hAD;
                    16'h6846: data_out = 8'hAE;
                    16'h6847: data_out = 8'hAF;
                    16'h6848: data_out = 8'hB0;
                    16'h6849: data_out = 8'hB1;
                    16'h684A: data_out = 8'hB2;
                    16'h684B: data_out = 8'hB3;
                    16'h684C: data_out = 8'hB4;
                    16'h684D: data_out = 8'hB5;
                    16'h684E: data_out = 8'hB6;
                    16'h684F: data_out = 8'hB7;
                    16'h6850: data_out = 8'hB8;
                    16'h6851: data_out = 8'hB9;
                    16'h6852: data_out = 8'hBA;
                    16'h6853: data_out = 8'hBB;
                    16'h6854: data_out = 8'hBC;
                    16'h6855: data_out = 8'hBD;
                    16'h6856: data_out = 8'hBE;
                    16'h6857: data_out = 8'hBF;
                    16'h6858: data_out = 8'hC0;
                    16'h6859: data_out = 8'hC1;
                    16'h685A: data_out = 8'hC2;
                    16'h685B: data_out = 8'hC3;
                    16'h685C: data_out = 8'hC4;
                    16'h685D: data_out = 8'hC5;
                    16'h685E: data_out = 8'hC6;
                    16'h685F: data_out = 8'hC7;
                    16'h6860: data_out = 8'hC8;
                    16'h6861: data_out = 8'hC9;
                    16'h6862: data_out = 8'hCA;
                    16'h6863: data_out = 8'hCB;
                    16'h6864: data_out = 8'hCC;
                    16'h6865: data_out = 8'hCD;
                    16'h6866: data_out = 8'hCE;
                    16'h6867: data_out = 8'hCF;
                    16'h6868: data_out = 8'hD0;
                    16'h6869: data_out = 8'hD1;
                    16'h686A: data_out = 8'hD2;
                    16'h686B: data_out = 8'hD3;
                    16'h686C: data_out = 8'hD4;
                    16'h686D: data_out = 8'hD5;
                    16'h686E: data_out = 8'hD6;
                    16'h686F: data_out = 8'hD7;
                    16'h6870: data_out = 8'hD8;
                    16'h6871: data_out = 8'hD9;
                    16'h6872: data_out = 8'hDA;
                    16'h6873: data_out = 8'hDB;
                    16'h6874: data_out = 8'hDC;
                    16'h6875: data_out = 8'hDD;
                    16'h6876: data_out = 8'hDE;
                    16'h6877: data_out = 8'hDF;
                    16'h6878: data_out = 8'hE0;
                    16'h6879: data_out = 8'hE1;
                    16'h687A: data_out = 8'hE2;
                    16'h687B: data_out = 8'hE3;
                    16'h687C: data_out = 8'hE4;
                    16'h687D: data_out = 8'hE5;
                    16'h687E: data_out = 8'hE6;
                    16'h687F: data_out = 8'hE7;
                    16'h6880: data_out = 8'h68;
                    16'h6881: data_out = 8'h67;
                    16'h6882: data_out = 8'h66;
                    16'h6883: data_out = 8'h65;
                    16'h6884: data_out = 8'h64;
                    16'h6885: data_out = 8'h63;
                    16'h6886: data_out = 8'h62;
                    16'h6887: data_out = 8'h61;
                    16'h6888: data_out = 8'h60;
                    16'h6889: data_out = 8'h5F;
                    16'h688A: data_out = 8'h5E;
                    16'h688B: data_out = 8'h5D;
                    16'h688C: data_out = 8'h5C;
                    16'h688D: data_out = 8'h5B;
                    16'h688E: data_out = 8'h5A;
                    16'h688F: data_out = 8'h59;
                    16'h6890: data_out = 8'h58;
                    16'h6891: data_out = 8'h57;
                    16'h6892: data_out = 8'h56;
                    16'h6893: data_out = 8'h55;
                    16'h6894: data_out = 8'h54;
                    16'h6895: data_out = 8'h53;
                    16'h6896: data_out = 8'h52;
                    16'h6897: data_out = 8'h51;
                    16'h6898: data_out = 8'h50;
                    16'h6899: data_out = 8'h4F;
                    16'h689A: data_out = 8'h4E;
                    16'h689B: data_out = 8'h4D;
                    16'h689C: data_out = 8'h4C;
                    16'h689D: data_out = 8'h4B;
                    16'h689E: data_out = 8'h4A;
                    16'h689F: data_out = 8'h49;
                    16'h68A0: data_out = 8'h48;
                    16'h68A1: data_out = 8'h47;
                    16'h68A2: data_out = 8'h46;
                    16'h68A3: data_out = 8'h45;
                    16'h68A4: data_out = 8'h44;
                    16'h68A5: data_out = 8'h43;
                    16'h68A6: data_out = 8'h42;
                    16'h68A7: data_out = 8'h41;
                    16'h68A8: data_out = 8'h40;
                    16'h68A9: data_out = 8'h3F;
                    16'h68AA: data_out = 8'h3E;
                    16'h68AB: data_out = 8'h3D;
                    16'h68AC: data_out = 8'h3C;
                    16'h68AD: data_out = 8'h3B;
                    16'h68AE: data_out = 8'h3A;
                    16'h68AF: data_out = 8'h39;
                    16'h68B0: data_out = 8'h38;
                    16'h68B1: data_out = 8'h37;
                    16'h68B2: data_out = 8'h36;
                    16'h68B3: data_out = 8'h35;
                    16'h68B4: data_out = 8'h34;
                    16'h68B5: data_out = 8'h33;
                    16'h68B6: data_out = 8'h32;
                    16'h68B7: data_out = 8'h31;
                    16'h68B8: data_out = 8'h30;
                    16'h68B9: data_out = 8'h2F;
                    16'h68BA: data_out = 8'h2E;
                    16'h68BB: data_out = 8'h2D;
                    16'h68BC: data_out = 8'h2C;
                    16'h68BD: data_out = 8'h2B;
                    16'h68BE: data_out = 8'h2A;
                    16'h68BF: data_out = 8'h29;
                    16'h68C0: data_out = 8'h28;
                    16'h68C1: data_out = 8'h27;
                    16'h68C2: data_out = 8'h26;
                    16'h68C3: data_out = 8'h25;
                    16'h68C4: data_out = 8'h24;
                    16'h68C5: data_out = 8'h23;
                    16'h68C6: data_out = 8'h22;
                    16'h68C7: data_out = 8'h21;
                    16'h68C8: data_out = 8'h20;
                    16'h68C9: data_out = 8'h1F;
                    16'h68CA: data_out = 8'h1E;
                    16'h68CB: data_out = 8'h1D;
                    16'h68CC: data_out = 8'h1C;
                    16'h68CD: data_out = 8'h1B;
                    16'h68CE: data_out = 8'h1A;
                    16'h68CF: data_out = 8'h19;
                    16'h68D0: data_out = 8'h18;
                    16'h68D1: data_out = 8'h17;
                    16'h68D2: data_out = 8'h16;
                    16'h68D3: data_out = 8'h15;
                    16'h68D4: data_out = 8'h14;
                    16'h68D5: data_out = 8'h13;
                    16'h68D6: data_out = 8'h12;
                    16'h68D7: data_out = 8'h11;
                    16'h68D8: data_out = 8'h10;
                    16'h68D9: data_out = 8'hF;
                    16'h68DA: data_out = 8'hE;
                    16'h68DB: data_out = 8'hD;
                    16'h68DC: data_out = 8'hC;
                    16'h68DD: data_out = 8'hB;
                    16'h68DE: data_out = 8'hA;
                    16'h68DF: data_out = 8'h9;
                    16'h68E0: data_out = 8'h8;
                    16'h68E1: data_out = 8'h7;
                    16'h68E2: data_out = 8'h6;
                    16'h68E3: data_out = 8'h5;
                    16'h68E4: data_out = 8'h4;
                    16'h68E5: data_out = 8'h3;
                    16'h68E6: data_out = 8'h2;
                    16'h68E7: data_out = 8'h1;
                    16'h68E8: data_out = 8'h0;
                    16'h68E9: data_out = 8'h81;
                    16'h68EA: data_out = 8'h82;
                    16'h68EB: data_out = 8'h83;
                    16'h68EC: data_out = 8'h84;
                    16'h68ED: data_out = 8'h85;
                    16'h68EE: data_out = 8'h86;
                    16'h68EF: data_out = 8'h87;
                    16'h68F0: data_out = 8'h88;
                    16'h68F1: data_out = 8'h89;
                    16'h68F2: data_out = 8'h8A;
                    16'h68F3: data_out = 8'h8B;
                    16'h68F4: data_out = 8'h8C;
                    16'h68F5: data_out = 8'h8D;
                    16'h68F6: data_out = 8'h8E;
                    16'h68F7: data_out = 8'h8F;
                    16'h68F8: data_out = 8'h90;
                    16'h68F9: data_out = 8'h91;
                    16'h68FA: data_out = 8'h92;
                    16'h68FB: data_out = 8'h93;
                    16'h68FC: data_out = 8'h94;
                    16'h68FD: data_out = 8'h95;
                    16'h68FE: data_out = 8'h96;
                    16'h68FF: data_out = 8'h97;
                    16'h6900: data_out = 8'h69;
                    16'h6901: data_out = 8'h6A;
                    16'h6902: data_out = 8'h6B;
                    16'h6903: data_out = 8'h6C;
                    16'h6904: data_out = 8'h6D;
                    16'h6905: data_out = 8'h6E;
                    16'h6906: data_out = 8'h6F;
                    16'h6907: data_out = 8'h70;
                    16'h6908: data_out = 8'h71;
                    16'h6909: data_out = 8'h72;
                    16'h690A: data_out = 8'h73;
                    16'h690B: data_out = 8'h74;
                    16'h690C: data_out = 8'h75;
                    16'h690D: data_out = 8'h76;
                    16'h690E: data_out = 8'h77;
                    16'h690F: data_out = 8'h78;
                    16'h6910: data_out = 8'h79;
                    16'h6911: data_out = 8'h7A;
                    16'h6912: data_out = 8'h7B;
                    16'h6913: data_out = 8'h7C;
                    16'h6914: data_out = 8'h7D;
                    16'h6915: data_out = 8'h7E;
                    16'h6916: data_out = 8'h7F;
                    16'h6917: data_out = 8'h80;
                    16'h6918: data_out = 8'h81;
                    16'h6919: data_out = 8'h82;
                    16'h691A: data_out = 8'h83;
                    16'h691B: data_out = 8'h84;
                    16'h691C: data_out = 8'h85;
                    16'h691D: data_out = 8'h86;
                    16'h691E: data_out = 8'h87;
                    16'h691F: data_out = 8'h88;
                    16'h6920: data_out = 8'h89;
                    16'h6921: data_out = 8'h8A;
                    16'h6922: data_out = 8'h8B;
                    16'h6923: data_out = 8'h8C;
                    16'h6924: data_out = 8'h8D;
                    16'h6925: data_out = 8'h8E;
                    16'h6926: data_out = 8'h8F;
                    16'h6927: data_out = 8'h90;
                    16'h6928: data_out = 8'h91;
                    16'h6929: data_out = 8'h92;
                    16'h692A: data_out = 8'h93;
                    16'h692B: data_out = 8'h94;
                    16'h692C: data_out = 8'h95;
                    16'h692D: data_out = 8'h96;
                    16'h692E: data_out = 8'h97;
                    16'h692F: data_out = 8'h98;
                    16'h6930: data_out = 8'h99;
                    16'h6931: data_out = 8'h9A;
                    16'h6932: data_out = 8'h9B;
                    16'h6933: data_out = 8'h9C;
                    16'h6934: data_out = 8'h9D;
                    16'h6935: data_out = 8'h9E;
                    16'h6936: data_out = 8'h9F;
                    16'h6937: data_out = 8'hA0;
                    16'h6938: data_out = 8'hA1;
                    16'h6939: data_out = 8'hA2;
                    16'h693A: data_out = 8'hA3;
                    16'h693B: data_out = 8'hA4;
                    16'h693C: data_out = 8'hA5;
                    16'h693D: data_out = 8'hA6;
                    16'h693E: data_out = 8'hA7;
                    16'h693F: data_out = 8'hA8;
                    16'h6940: data_out = 8'hA9;
                    16'h6941: data_out = 8'hAA;
                    16'h6942: data_out = 8'hAB;
                    16'h6943: data_out = 8'hAC;
                    16'h6944: data_out = 8'hAD;
                    16'h6945: data_out = 8'hAE;
                    16'h6946: data_out = 8'hAF;
                    16'h6947: data_out = 8'hB0;
                    16'h6948: data_out = 8'hB1;
                    16'h6949: data_out = 8'hB2;
                    16'h694A: data_out = 8'hB3;
                    16'h694B: data_out = 8'hB4;
                    16'h694C: data_out = 8'hB5;
                    16'h694D: data_out = 8'hB6;
                    16'h694E: data_out = 8'hB7;
                    16'h694F: data_out = 8'hB8;
                    16'h6950: data_out = 8'hB9;
                    16'h6951: data_out = 8'hBA;
                    16'h6952: data_out = 8'hBB;
                    16'h6953: data_out = 8'hBC;
                    16'h6954: data_out = 8'hBD;
                    16'h6955: data_out = 8'hBE;
                    16'h6956: data_out = 8'hBF;
                    16'h6957: data_out = 8'hC0;
                    16'h6958: data_out = 8'hC1;
                    16'h6959: data_out = 8'hC2;
                    16'h695A: data_out = 8'hC3;
                    16'h695B: data_out = 8'hC4;
                    16'h695C: data_out = 8'hC5;
                    16'h695D: data_out = 8'hC6;
                    16'h695E: data_out = 8'hC7;
                    16'h695F: data_out = 8'hC8;
                    16'h6960: data_out = 8'hC9;
                    16'h6961: data_out = 8'hCA;
                    16'h6962: data_out = 8'hCB;
                    16'h6963: data_out = 8'hCC;
                    16'h6964: data_out = 8'hCD;
                    16'h6965: data_out = 8'hCE;
                    16'h6966: data_out = 8'hCF;
                    16'h6967: data_out = 8'hD0;
                    16'h6968: data_out = 8'hD1;
                    16'h6969: data_out = 8'hD2;
                    16'h696A: data_out = 8'hD3;
                    16'h696B: data_out = 8'hD4;
                    16'h696C: data_out = 8'hD5;
                    16'h696D: data_out = 8'hD6;
                    16'h696E: data_out = 8'hD7;
                    16'h696F: data_out = 8'hD8;
                    16'h6970: data_out = 8'hD9;
                    16'h6971: data_out = 8'hDA;
                    16'h6972: data_out = 8'hDB;
                    16'h6973: data_out = 8'hDC;
                    16'h6974: data_out = 8'hDD;
                    16'h6975: data_out = 8'hDE;
                    16'h6976: data_out = 8'hDF;
                    16'h6977: data_out = 8'hE0;
                    16'h6978: data_out = 8'hE1;
                    16'h6979: data_out = 8'hE2;
                    16'h697A: data_out = 8'hE3;
                    16'h697B: data_out = 8'hE4;
                    16'h697C: data_out = 8'hE5;
                    16'h697D: data_out = 8'hE6;
                    16'h697E: data_out = 8'hE7;
                    16'h697F: data_out = 8'hE8;
                    16'h6980: data_out = 8'h69;
                    16'h6981: data_out = 8'h68;
                    16'h6982: data_out = 8'h67;
                    16'h6983: data_out = 8'h66;
                    16'h6984: data_out = 8'h65;
                    16'h6985: data_out = 8'h64;
                    16'h6986: data_out = 8'h63;
                    16'h6987: data_out = 8'h62;
                    16'h6988: data_out = 8'h61;
                    16'h6989: data_out = 8'h60;
                    16'h698A: data_out = 8'h5F;
                    16'h698B: data_out = 8'h5E;
                    16'h698C: data_out = 8'h5D;
                    16'h698D: data_out = 8'h5C;
                    16'h698E: data_out = 8'h5B;
                    16'h698F: data_out = 8'h5A;
                    16'h6990: data_out = 8'h59;
                    16'h6991: data_out = 8'h58;
                    16'h6992: data_out = 8'h57;
                    16'h6993: data_out = 8'h56;
                    16'h6994: data_out = 8'h55;
                    16'h6995: data_out = 8'h54;
                    16'h6996: data_out = 8'h53;
                    16'h6997: data_out = 8'h52;
                    16'h6998: data_out = 8'h51;
                    16'h6999: data_out = 8'h50;
                    16'h699A: data_out = 8'h4F;
                    16'h699B: data_out = 8'h4E;
                    16'h699C: data_out = 8'h4D;
                    16'h699D: data_out = 8'h4C;
                    16'h699E: data_out = 8'h4B;
                    16'h699F: data_out = 8'h4A;
                    16'h69A0: data_out = 8'h49;
                    16'h69A1: data_out = 8'h48;
                    16'h69A2: data_out = 8'h47;
                    16'h69A3: data_out = 8'h46;
                    16'h69A4: data_out = 8'h45;
                    16'h69A5: data_out = 8'h44;
                    16'h69A6: data_out = 8'h43;
                    16'h69A7: data_out = 8'h42;
                    16'h69A8: data_out = 8'h41;
                    16'h69A9: data_out = 8'h40;
                    16'h69AA: data_out = 8'h3F;
                    16'h69AB: data_out = 8'h3E;
                    16'h69AC: data_out = 8'h3D;
                    16'h69AD: data_out = 8'h3C;
                    16'h69AE: data_out = 8'h3B;
                    16'h69AF: data_out = 8'h3A;
                    16'h69B0: data_out = 8'h39;
                    16'h69B1: data_out = 8'h38;
                    16'h69B2: data_out = 8'h37;
                    16'h69B3: data_out = 8'h36;
                    16'h69B4: data_out = 8'h35;
                    16'h69B5: data_out = 8'h34;
                    16'h69B6: data_out = 8'h33;
                    16'h69B7: data_out = 8'h32;
                    16'h69B8: data_out = 8'h31;
                    16'h69B9: data_out = 8'h30;
                    16'h69BA: data_out = 8'h2F;
                    16'h69BB: data_out = 8'h2E;
                    16'h69BC: data_out = 8'h2D;
                    16'h69BD: data_out = 8'h2C;
                    16'h69BE: data_out = 8'h2B;
                    16'h69BF: data_out = 8'h2A;
                    16'h69C0: data_out = 8'h29;
                    16'h69C1: data_out = 8'h28;
                    16'h69C2: data_out = 8'h27;
                    16'h69C3: data_out = 8'h26;
                    16'h69C4: data_out = 8'h25;
                    16'h69C5: data_out = 8'h24;
                    16'h69C6: data_out = 8'h23;
                    16'h69C7: data_out = 8'h22;
                    16'h69C8: data_out = 8'h21;
                    16'h69C9: data_out = 8'h20;
                    16'h69CA: data_out = 8'h1F;
                    16'h69CB: data_out = 8'h1E;
                    16'h69CC: data_out = 8'h1D;
                    16'h69CD: data_out = 8'h1C;
                    16'h69CE: data_out = 8'h1B;
                    16'h69CF: data_out = 8'h1A;
                    16'h69D0: data_out = 8'h19;
                    16'h69D1: data_out = 8'h18;
                    16'h69D2: data_out = 8'h17;
                    16'h69D3: data_out = 8'h16;
                    16'h69D4: data_out = 8'h15;
                    16'h69D5: data_out = 8'h14;
                    16'h69D6: data_out = 8'h13;
                    16'h69D7: data_out = 8'h12;
                    16'h69D8: data_out = 8'h11;
                    16'h69D9: data_out = 8'h10;
                    16'h69DA: data_out = 8'hF;
                    16'h69DB: data_out = 8'hE;
                    16'h69DC: data_out = 8'hD;
                    16'h69DD: data_out = 8'hC;
                    16'h69DE: data_out = 8'hB;
                    16'h69DF: data_out = 8'hA;
                    16'h69E0: data_out = 8'h9;
                    16'h69E1: data_out = 8'h8;
                    16'h69E2: data_out = 8'h7;
                    16'h69E3: data_out = 8'h6;
                    16'h69E4: data_out = 8'h5;
                    16'h69E5: data_out = 8'h4;
                    16'h69E6: data_out = 8'h3;
                    16'h69E7: data_out = 8'h2;
                    16'h69E8: data_out = 8'h1;
                    16'h69E9: data_out = 8'h0;
                    16'h69EA: data_out = 8'h81;
                    16'h69EB: data_out = 8'h82;
                    16'h69EC: data_out = 8'h83;
                    16'h69ED: data_out = 8'h84;
                    16'h69EE: data_out = 8'h85;
                    16'h69EF: data_out = 8'h86;
                    16'h69F0: data_out = 8'h87;
                    16'h69F1: data_out = 8'h88;
                    16'h69F2: data_out = 8'h89;
                    16'h69F3: data_out = 8'h8A;
                    16'h69F4: data_out = 8'h8B;
                    16'h69F5: data_out = 8'h8C;
                    16'h69F6: data_out = 8'h8D;
                    16'h69F7: data_out = 8'h8E;
                    16'h69F8: data_out = 8'h8F;
                    16'h69F9: data_out = 8'h90;
                    16'h69FA: data_out = 8'h91;
                    16'h69FB: data_out = 8'h92;
                    16'h69FC: data_out = 8'h93;
                    16'h69FD: data_out = 8'h94;
                    16'h69FE: data_out = 8'h95;
                    16'h69FF: data_out = 8'h96;
                    16'h6A00: data_out = 8'h6A;
                    16'h6A01: data_out = 8'h6B;
                    16'h6A02: data_out = 8'h6C;
                    16'h6A03: data_out = 8'h6D;
                    16'h6A04: data_out = 8'h6E;
                    16'h6A05: data_out = 8'h6F;
                    16'h6A06: data_out = 8'h70;
                    16'h6A07: data_out = 8'h71;
                    16'h6A08: data_out = 8'h72;
                    16'h6A09: data_out = 8'h73;
                    16'h6A0A: data_out = 8'h74;
                    16'h6A0B: data_out = 8'h75;
                    16'h6A0C: data_out = 8'h76;
                    16'h6A0D: data_out = 8'h77;
                    16'h6A0E: data_out = 8'h78;
                    16'h6A0F: data_out = 8'h79;
                    16'h6A10: data_out = 8'h7A;
                    16'h6A11: data_out = 8'h7B;
                    16'h6A12: data_out = 8'h7C;
                    16'h6A13: data_out = 8'h7D;
                    16'h6A14: data_out = 8'h7E;
                    16'h6A15: data_out = 8'h7F;
                    16'h6A16: data_out = 8'h80;
                    16'h6A17: data_out = 8'h81;
                    16'h6A18: data_out = 8'h82;
                    16'h6A19: data_out = 8'h83;
                    16'h6A1A: data_out = 8'h84;
                    16'h6A1B: data_out = 8'h85;
                    16'h6A1C: data_out = 8'h86;
                    16'h6A1D: data_out = 8'h87;
                    16'h6A1E: data_out = 8'h88;
                    16'h6A1F: data_out = 8'h89;
                    16'h6A20: data_out = 8'h8A;
                    16'h6A21: data_out = 8'h8B;
                    16'h6A22: data_out = 8'h8C;
                    16'h6A23: data_out = 8'h8D;
                    16'h6A24: data_out = 8'h8E;
                    16'h6A25: data_out = 8'h8F;
                    16'h6A26: data_out = 8'h90;
                    16'h6A27: data_out = 8'h91;
                    16'h6A28: data_out = 8'h92;
                    16'h6A29: data_out = 8'h93;
                    16'h6A2A: data_out = 8'h94;
                    16'h6A2B: data_out = 8'h95;
                    16'h6A2C: data_out = 8'h96;
                    16'h6A2D: data_out = 8'h97;
                    16'h6A2E: data_out = 8'h98;
                    16'h6A2F: data_out = 8'h99;
                    16'h6A30: data_out = 8'h9A;
                    16'h6A31: data_out = 8'h9B;
                    16'h6A32: data_out = 8'h9C;
                    16'h6A33: data_out = 8'h9D;
                    16'h6A34: data_out = 8'h9E;
                    16'h6A35: data_out = 8'h9F;
                    16'h6A36: data_out = 8'hA0;
                    16'h6A37: data_out = 8'hA1;
                    16'h6A38: data_out = 8'hA2;
                    16'h6A39: data_out = 8'hA3;
                    16'h6A3A: data_out = 8'hA4;
                    16'h6A3B: data_out = 8'hA5;
                    16'h6A3C: data_out = 8'hA6;
                    16'h6A3D: data_out = 8'hA7;
                    16'h6A3E: data_out = 8'hA8;
                    16'h6A3F: data_out = 8'hA9;
                    16'h6A40: data_out = 8'hAA;
                    16'h6A41: data_out = 8'hAB;
                    16'h6A42: data_out = 8'hAC;
                    16'h6A43: data_out = 8'hAD;
                    16'h6A44: data_out = 8'hAE;
                    16'h6A45: data_out = 8'hAF;
                    16'h6A46: data_out = 8'hB0;
                    16'h6A47: data_out = 8'hB1;
                    16'h6A48: data_out = 8'hB2;
                    16'h6A49: data_out = 8'hB3;
                    16'h6A4A: data_out = 8'hB4;
                    16'h6A4B: data_out = 8'hB5;
                    16'h6A4C: data_out = 8'hB6;
                    16'h6A4D: data_out = 8'hB7;
                    16'h6A4E: data_out = 8'hB8;
                    16'h6A4F: data_out = 8'hB9;
                    16'h6A50: data_out = 8'hBA;
                    16'h6A51: data_out = 8'hBB;
                    16'h6A52: data_out = 8'hBC;
                    16'h6A53: data_out = 8'hBD;
                    16'h6A54: data_out = 8'hBE;
                    16'h6A55: data_out = 8'hBF;
                    16'h6A56: data_out = 8'hC0;
                    16'h6A57: data_out = 8'hC1;
                    16'h6A58: data_out = 8'hC2;
                    16'h6A59: data_out = 8'hC3;
                    16'h6A5A: data_out = 8'hC4;
                    16'h6A5B: data_out = 8'hC5;
                    16'h6A5C: data_out = 8'hC6;
                    16'h6A5D: data_out = 8'hC7;
                    16'h6A5E: data_out = 8'hC8;
                    16'h6A5F: data_out = 8'hC9;
                    16'h6A60: data_out = 8'hCA;
                    16'h6A61: data_out = 8'hCB;
                    16'h6A62: data_out = 8'hCC;
                    16'h6A63: data_out = 8'hCD;
                    16'h6A64: data_out = 8'hCE;
                    16'h6A65: data_out = 8'hCF;
                    16'h6A66: data_out = 8'hD0;
                    16'h6A67: data_out = 8'hD1;
                    16'h6A68: data_out = 8'hD2;
                    16'h6A69: data_out = 8'hD3;
                    16'h6A6A: data_out = 8'hD4;
                    16'h6A6B: data_out = 8'hD5;
                    16'h6A6C: data_out = 8'hD6;
                    16'h6A6D: data_out = 8'hD7;
                    16'h6A6E: data_out = 8'hD8;
                    16'h6A6F: data_out = 8'hD9;
                    16'h6A70: data_out = 8'hDA;
                    16'h6A71: data_out = 8'hDB;
                    16'h6A72: data_out = 8'hDC;
                    16'h6A73: data_out = 8'hDD;
                    16'h6A74: data_out = 8'hDE;
                    16'h6A75: data_out = 8'hDF;
                    16'h6A76: data_out = 8'hE0;
                    16'h6A77: data_out = 8'hE1;
                    16'h6A78: data_out = 8'hE2;
                    16'h6A79: data_out = 8'hE3;
                    16'h6A7A: data_out = 8'hE4;
                    16'h6A7B: data_out = 8'hE5;
                    16'h6A7C: data_out = 8'hE6;
                    16'h6A7D: data_out = 8'hE7;
                    16'h6A7E: data_out = 8'hE8;
                    16'h6A7F: data_out = 8'hE9;
                    16'h6A80: data_out = 8'h6A;
                    16'h6A81: data_out = 8'h69;
                    16'h6A82: data_out = 8'h68;
                    16'h6A83: data_out = 8'h67;
                    16'h6A84: data_out = 8'h66;
                    16'h6A85: data_out = 8'h65;
                    16'h6A86: data_out = 8'h64;
                    16'h6A87: data_out = 8'h63;
                    16'h6A88: data_out = 8'h62;
                    16'h6A89: data_out = 8'h61;
                    16'h6A8A: data_out = 8'h60;
                    16'h6A8B: data_out = 8'h5F;
                    16'h6A8C: data_out = 8'h5E;
                    16'h6A8D: data_out = 8'h5D;
                    16'h6A8E: data_out = 8'h5C;
                    16'h6A8F: data_out = 8'h5B;
                    16'h6A90: data_out = 8'h5A;
                    16'h6A91: data_out = 8'h59;
                    16'h6A92: data_out = 8'h58;
                    16'h6A93: data_out = 8'h57;
                    16'h6A94: data_out = 8'h56;
                    16'h6A95: data_out = 8'h55;
                    16'h6A96: data_out = 8'h54;
                    16'h6A97: data_out = 8'h53;
                    16'h6A98: data_out = 8'h52;
                    16'h6A99: data_out = 8'h51;
                    16'h6A9A: data_out = 8'h50;
                    16'h6A9B: data_out = 8'h4F;
                    16'h6A9C: data_out = 8'h4E;
                    16'h6A9D: data_out = 8'h4D;
                    16'h6A9E: data_out = 8'h4C;
                    16'h6A9F: data_out = 8'h4B;
                    16'h6AA0: data_out = 8'h4A;
                    16'h6AA1: data_out = 8'h49;
                    16'h6AA2: data_out = 8'h48;
                    16'h6AA3: data_out = 8'h47;
                    16'h6AA4: data_out = 8'h46;
                    16'h6AA5: data_out = 8'h45;
                    16'h6AA6: data_out = 8'h44;
                    16'h6AA7: data_out = 8'h43;
                    16'h6AA8: data_out = 8'h42;
                    16'h6AA9: data_out = 8'h41;
                    16'h6AAA: data_out = 8'h40;
                    16'h6AAB: data_out = 8'h3F;
                    16'h6AAC: data_out = 8'h3E;
                    16'h6AAD: data_out = 8'h3D;
                    16'h6AAE: data_out = 8'h3C;
                    16'h6AAF: data_out = 8'h3B;
                    16'h6AB0: data_out = 8'h3A;
                    16'h6AB1: data_out = 8'h39;
                    16'h6AB2: data_out = 8'h38;
                    16'h6AB3: data_out = 8'h37;
                    16'h6AB4: data_out = 8'h36;
                    16'h6AB5: data_out = 8'h35;
                    16'h6AB6: data_out = 8'h34;
                    16'h6AB7: data_out = 8'h33;
                    16'h6AB8: data_out = 8'h32;
                    16'h6AB9: data_out = 8'h31;
                    16'h6ABA: data_out = 8'h30;
                    16'h6ABB: data_out = 8'h2F;
                    16'h6ABC: data_out = 8'h2E;
                    16'h6ABD: data_out = 8'h2D;
                    16'h6ABE: data_out = 8'h2C;
                    16'h6ABF: data_out = 8'h2B;
                    16'h6AC0: data_out = 8'h2A;
                    16'h6AC1: data_out = 8'h29;
                    16'h6AC2: data_out = 8'h28;
                    16'h6AC3: data_out = 8'h27;
                    16'h6AC4: data_out = 8'h26;
                    16'h6AC5: data_out = 8'h25;
                    16'h6AC6: data_out = 8'h24;
                    16'h6AC7: data_out = 8'h23;
                    16'h6AC8: data_out = 8'h22;
                    16'h6AC9: data_out = 8'h21;
                    16'h6ACA: data_out = 8'h20;
                    16'h6ACB: data_out = 8'h1F;
                    16'h6ACC: data_out = 8'h1E;
                    16'h6ACD: data_out = 8'h1D;
                    16'h6ACE: data_out = 8'h1C;
                    16'h6ACF: data_out = 8'h1B;
                    16'h6AD0: data_out = 8'h1A;
                    16'h6AD1: data_out = 8'h19;
                    16'h6AD2: data_out = 8'h18;
                    16'h6AD3: data_out = 8'h17;
                    16'h6AD4: data_out = 8'h16;
                    16'h6AD5: data_out = 8'h15;
                    16'h6AD6: data_out = 8'h14;
                    16'h6AD7: data_out = 8'h13;
                    16'h6AD8: data_out = 8'h12;
                    16'h6AD9: data_out = 8'h11;
                    16'h6ADA: data_out = 8'h10;
                    16'h6ADB: data_out = 8'hF;
                    16'h6ADC: data_out = 8'hE;
                    16'h6ADD: data_out = 8'hD;
                    16'h6ADE: data_out = 8'hC;
                    16'h6ADF: data_out = 8'hB;
                    16'h6AE0: data_out = 8'hA;
                    16'h6AE1: data_out = 8'h9;
                    16'h6AE2: data_out = 8'h8;
                    16'h6AE3: data_out = 8'h7;
                    16'h6AE4: data_out = 8'h6;
                    16'h6AE5: data_out = 8'h5;
                    16'h6AE6: data_out = 8'h4;
                    16'h6AE7: data_out = 8'h3;
                    16'h6AE8: data_out = 8'h2;
                    16'h6AE9: data_out = 8'h1;
                    16'h6AEA: data_out = 8'h0;
                    16'h6AEB: data_out = 8'h81;
                    16'h6AEC: data_out = 8'h82;
                    16'h6AED: data_out = 8'h83;
                    16'h6AEE: data_out = 8'h84;
                    16'h6AEF: data_out = 8'h85;
                    16'h6AF0: data_out = 8'h86;
                    16'h6AF1: data_out = 8'h87;
                    16'h6AF2: data_out = 8'h88;
                    16'h6AF3: data_out = 8'h89;
                    16'h6AF4: data_out = 8'h8A;
                    16'h6AF5: data_out = 8'h8B;
                    16'h6AF6: data_out = 8'h8C;
                    16'h6AF7: data_out = 8'h8D;
                    16'h6AF8: data_out = 8'h8E;
                    16'h6AF9: data_out = 8'h8F;
                    16'h6AFA: data_out = 8'h90;
                    16'h6AFB: data_out = 8'h91;
                    16'h6AFC: data_out = 8'h92;
                    16'h6AFD: data_out = 8'h93;
                    16'h6AFE: data_out = 8'h94;
                    16'h6AFF: data_out = 8'h95;
                    16'h6B00: data_out = 8'h6B;
                    16'h6B01: data_out = 8'h6C;
                    16'h6B02: data_out = 8'h6D;
                    16'h6B03: data_out = 8'h6E;
                    16'h6B04: data_out = 8'h6F;
                    16'h6B05: data_out = 8'h70;
                    16'h6B06: data_out = 8'h71;
                    16'h6B07: data_out = 8'h72;
                    16'h6B08: data_out = 8'h73;
                    16'h6B09: data_out = 8'h74;
                    16'h6B0A: data_out = 8'h75;
                    16'h6B0B: data_out = 8'h76;
                    16'h6B0C: data_out = 8'h77;
                    16'h6B0D: data_out = 8'h78;
                    16'h6B0E: data_out = 8'h79;
                    16'h6B0F: data_out = 8'h7A;
                    16'h6B10: data_out = 8'h7B;
                    16'h6B11: data_out = 8'h7C;
                    16'h6B12: data_out = 8'h7D;
                    16'h6B13: data_out = 8'h7E;
                    16'h6B14: data_out = 8'h7F;
                    16'h6B15: data_out = 8'h80;
                    16'h6B16: data_out = 8'h81;
                    16'h6B17: data_out = 8'h82;
                    16'h6B18: data_out = 8'h83;
                    16'h6B19: data_out = 8'h84;
                    16'h6B1A: data_out = 8'h85;
                    16'h6B1B: data_out = 8'h86;
                    16'h6B1C: data_out = 8'h87;
                    16'h6B1D: data_out = 8'h88;
                    16'h6B1E: data_out = 8'h89;
                    16'h6B1F: data_out = 8'h8A;
                    16'h6B20: data_out = 8'h8B;
                    16'h6B21: data_out = 8'h8C;
                    16'h6B22: data_out = 8'h8D;
                    16'h6B23: data_out = 8'h8E;
                    16'h6B24: data_out = 8'h8F;
                    16'h6B25: data_out = 8'h90;
                    16'h6B26: data_out = 8'h91;
                    16'h6B27: data_out = 8'h92;
                    16'h6B28: data_out = 8'h93;
                    16'h6B29: data_out = 8'h94;
                    16'h6B2A: data_out = 8'h95;
                    16'h6B2B: data_out = 8'h96;
                    16'h6B2C: data_out = 8'h97;
                    16'h6B2D: data_out = 8'h98;
                    16'h6B2E: data_out = 8'h99;
                    16'h6B2F: data_out = 8'h9A;
                    16'h6B30: data_out = 8'h9B;
                    16'h6B31: data_out = 8'h9C;
                    16'h6B32: data_out = 8'h9D;
                    16'h6B33: data_out = 8'h9E;
                    16'h6B34: data_out = 8'h9F;
                    16'h6B35: data_out = 8'hA0;
                    16'h6B36: data_out = 8'hA1;
                    16'h6B37: data_out = 8'hA2;
                    16'h6B38: data_out = 8'hA3;
                    16'h6B39: data_out = 8'hA4;
                    16'h6B3A: data_out = 8'hA5;
                    16'h6B3B: data_out = 8'hA6;
                    16'h6B3C: data_out = 8'hA7;
                    16'h6B3D: data_out = 8'hA8;
                    16'h6B3E: data_out = 8'hA9;
                    16'h6B3F: data_out = 8'hAA;
                    16'h6B40: data_out = 8'hAB;
                    16'h6B41: data_out = 8'hAC;
                    16'h6B42: data_out = 8'hAD;
                    16'h6B43: data_out = 8'hAE;
                    16'h6B44: data_out = 8'hAF;
                    16'h6B45: data_out = 8'hB0;
                    16'h6B46: data_out = 8'hB1;
                    16'h6B47: data_out = 8'hB2;
                    16'h6B48: data_out = 8'hB3;
                    16'h6B49: data_out = 8'hB4;
                    16'h6B4A: data_out = 8'hB5;
                    16'h6B4B: data_out = 8'hB6;
                    16'h6B4C: data_out = 8'hB7;
                    16'h6B4D: data_out = 8'hB8;
                    16'h6B4E: data_out = 8'hB9;
                    16'h6B4F: data_out = 8'hBA;
                    16'h6B50: data_out = 8'hBB;
                    16'h6B51: data_out = 8'hBC;
                    16'h6B52: data_out = 8'hBD;
                    16'h6B53: data_out = 8'hBE;
                    16'h6B54: data_out = 8'hBF;
                    16'h6B55: data_out = 8'hC0;
                    16'h6B56: data_out = 8'hC1;
                    16'h6B57: data_out = 8'hC2;
                    16'h6B58: data_out = 8'hC3;
                    16'h6B59: data_out = 8'hC4;
                    16'h6B5A: data_out = 8'hC5;
                    16'h6B5B: data_out = 8'hC6;
                    16'h6B5C: data_out = 8'hC7;
                    16'h6B5D: data_out = 8'hC8;
                    16'h6B5E: data_out = 8'hC9;
                    16'h6B5F: data_out = 8'hCA;
                    16'h6B60: data_out = 8'hCB;
                    16'h6B61: data_out = 8'hCC;
                    16'h6B62: data_out = 8'hCD;
                    16'h6B63: data_out = 8'hCE;
                    16'h6B64: data_out = 8'hCF;
                    16'h6B65: data_out = 8'hD0;
                    16'h6B66: data_out = 8'hD1;
                    16'h6B67: data_out = 8'hD2;
                    16'h6B68: data_out = 8'hD3;
                    16'h6B69: data_out = 8'hD4;
                    16'h6B6A: data_out = 8'hD5;
                    16'h6B6B: data_out = 8'hD6;
                    16'h6B6C: data_out = 8'hD7;
                    16'h6B6D: data_out = 8'hD8;
                    16'h6B6E: data_out = 8'hD9;
                    16'h6B6F: data_out = 8'hDA;
                    16'h6B70: data_out = 8'hDB;
                    16'h6B71: data_out = 8'hDC;
                    16'h6B72: data_out = 8'hDD;
                    16'h6B73: data_out = 8'hDE;
                    16'h6B74: data_out = 8'hDF;
                    16'h6B75: data_out = 8'hE0;
                    16'h6B76: data_out = 8'hE1;
                    16'h6B77: data_out = 8'hE2;
                    16'h6B78: data_out = 8'hE3;
                    16'h6B79: data_out = 8'hE4;
                    16'h6B7A: data_out = 8'hE5;
                    16'h6B7B: data_out = 8'hE6;
                    16'h6B7C: data_out = 8'hE7;
                    16'h6B7D: data_out = 8'hE8;
                    16'h6B7E: data_out = 8'hE9;
                    16'h6B7F: data_out = 8'hEA;
                    16'h6B80: data_out = 8'h6B;
                    16'h6B81: data_out = 8'h6A;
                    16'h6B82: data_out = 8'h69;
                    16'h6B83: data_out = 8'h68;
                    16'h6B84: data_out = 8'h67;
                    16'h6B85: data_out = 8'h66;
                    16'h6B86: data_out = 8'h65;
                    16'h6B87: data_out = 8'h64;
                    16'h6B88: data_out = 8'h63;
                    16'h6B89: data_out = 8'h62;
                    16'h6B8A: data_out = 8'h61;
                    16'h6B8B: data_out = 8'h60;
                    16'h6B8C: data_out = 8'h5F;
                    16'h6B8D: data_out = 8'h5E;
                    16'h6B8E: data_out = 8'h5D;
                    16'h6B8F: data_out = 8'h5C;
                    16'h6B90: data_out = 8'h5B;
                    16'h6B91: data_out = 8'h5A;
                    16'h6B92: data_out = 8'h59;
                    16'h6B93: data_out = 8'h58;
                    16'h6B94: data_out = 8'h57;
                    16'h6B95: data_out = 8'h56;
                    16'h6B96: data_out = 8'h55;
                    16'h6B97: data_out = 8'h54;
                    16'h6B98: data_out = 8'h53;
                    16'h6B99: data_out = 8'h52;
                    16'h6B9A: data_out = 8'h51;
                    16'h6B9B: data_out = 8'h50;
                    16'h6B9C: data_out = 8'h4F;
                    16'h6B9D: data_out = 8'h4E;
                    16'h6B9E: data_out = 8'h4D;
                    16'h6B9F: data_out = 8'h4C;
                    16'h6BA0: data_out = 8'h4B;
                    16'h6BA1: data_out = 8'h4A;
                    16'h6BA2: data_out = 8'h49;
                    16'h6BA3: data_out = 8'h48;
                    16'h6BA4: data_out = 8'h47;
                    16'h6BA5: data_out = 8'h46;
                    16'h6BA6: data_out = 8'h45;
                    16'h6BA7: data_out = 8'h44;
                    16'h6BA8: data_out = 8'h43;
                    16'h6BA9: data_out = 8'h42;
                    16'h6BAA: data_out = 8'h41;
                    16'h6BAB: data_out = 8'h40;
                    16'h6BAC: data_out = 8'h3F;
                    16'h6BAD: data_out = 8'h3E;
                    16'h6BAE: data_out = 8'h3D;
                    16'h6BAF: data_out = 8'h3C;
                    16'h6BB0: data_out = 8'h3B;
                    16'h6BB1: data_out = 8'h3A;
                    16'h6BB2: data_out = 8'h39;
                    16'h6BB3: data_out = 8'h38;
                    16'h6BB4: data_out = 8'h37;
                    16'h6BB5: data_out = 8'h36;
                    16'h6BB6: data_out = 8'h35;
                    16'h6BB7: data_out = 8'h34;
                    16'h6BB8: data_out = 8'h33;
                    16'h6BB9: data_out = 8'h32;
                    16'h6BBA: data_out = 8'h31;
                    16'h6BBB: data_out = 8'h30;
                    16'h6BBC: data_out = 8'h2F;
                    16'h6BBD: data_out = 8'h2E;
                    16'h6BBE: data_out = 8'h2D;
                    16'h6BBF: data_out = 8'h2C;
                    16'h6BC0: data_out = 8'h2B;
                    16'h6BC1: data_out = 8'h2A;
                    16'h6BC2: data_out = 8'h29;
                    16'h6BC3: data_out = 8'h28;
                    16'h6BC4: data_out = 8'h27;
                    16'h6BC5: data_out = 8'h26;
                    16'h6BC6: data_out = 8'h25;
                    16'h6BC7: data_out = 8'h24;
                    16'h6BC8: data_out = 8'h23;
                    16'h6BC9: data_out = 8'h22;
                    16'h6BCA: data_out = 8'h21;
                    16'h6BCB: data_out = 8'h20;
                    16'h6BCC: data_out = 8'h1F;
                    16'h6BCD: data_out = 8'h1E;
                    16'h6BCE: data_out = 8'h1D;
                    16'h6BCF: data_out = 8'h1C;
                    16'h6BD0: data_out = 8'h1B;
                    16'h6BD1: data_out = 8'h1A;
                    16'h6BD2: data_out = 8'h19;
                    16'h6BD3: data_out = 8'h18;
                    16'h6BD4: data_out = 8'h17;
                    16'h6BD5: data_out = 8'h16;
                    16'h6BD6: data_out = 8'h15;
                    16'h6BD7: data_out = 8'h14;
                    16'h6BD8: data_out = 8'h13;
                    16'h6BD9: data_out = 8'h12;
                    16'h6BDA: data_out = 8'h11;
                    16'h6BDB: data_out = 8'h10;
                    16'h6BDC: data_out = 8'hF;
                    16'h6BDD: data_out = 8'hE;
                    16'h6BDE: data_out = 8'hD;
                    16'h6BDF: data_out = 8'hC;
                    16'h6BE0: data_out = 8'hB;
                    16'h6BE1: data_out = 8'hA;
                    16'h6BE2: data_out = 8'h9;
                    16'h6BE3: data_out = 8'h8;
                    16'h6BE4: data_out = 8'h7;
                    16'h6BE5: data_out = 8'h6;
                    16'h6BE6: data_out = 8'h5;
                    16'h6BE7: data_out = 8'h4;
                    16'h6BE8: data_out = 8'h3;
                    16'h6BE9: data_out = 8'h2;
                    16'h6BEA: data_out = 8'h1;
                    16'h6BEB: data_out = 8'h0;
                    16'h6BEC: data_out = 8'h81;
                    16'h6BED: data_out = 8'h82;
                    16'h6BEE: data_out = 8'h83;
                    16'h6BEF: data_out = 8'h84;
                    16'h6BF0: data_out = 8'h85;
                    16'h6BF1: data_out = 8'h86;
                    16'h6BF2: data_out = 8'h87;
                    16'h6BF3: data_out = 8'h88;
                    16'h6BF4: data_out = 8'h89;
                    16'h6BF5: data_out = 8'h8A;
                    16'h6BF6: data_out = 8'h8B;
                    16'h6BF7: data_out = 8'h8C;
                    16'h6BF8: data_out = 8'h8D;
                    16'h6BF9: data_out = 8'h8E;
                    16'h6BFA: data_out = 8'h8F;
                    16'h6BFB: data_out = 8'h90;
                    16'h6BFC: data_out = 8'h91;
                    16'h6BFD: data_out = 8'h92;
                    16'h6BFE: data_out = 8'h93;
                    16'h6BFF: data_out = 8'h94;
                    16'h6C00: data_out = 8'h6C;
                    16'h6C01: data_out = 8'h6D;
                    16'h6C02: data_out = 8'h6E;
                    16'h6C03: data_out = 8'h6F;
                    16'h6C04: data_out = 8'h70;
                    16'h6C05: data_out = 8'h71;
                    16'h6C06: data_out = 8'h72;
                    16'h6C07: data_out = 8'h73;
                    16'h6C08: data_out = 8'h74;
                    16'h6C09: data_out = 8'h75;
                    16'h6C0A: data_out = 8'h76;
                    16'h6C0B: data_out = 8'h77;
                    16'h6C0C: data_out = 8'h78;
                    16'h6C0D: data_out = 8'h79;
                    16'h6C0E: data_out = 8'h7A;
                    16'h6C0F: data_out = 8'h7B;
                    16'h6C10: data_out = 8'h7C;
                    16'h6C11: data_out = 8'h7D;
                    16'h6C12: data_out = 8'h7E;
                    16'h6C13: data_out = 8'h7F;
                    16'h6C14: data_out = 8'h80;
                    16'h6C15: data_out = 8'h81;
                    16'h6C16: data_out = 8'h82;
                    16'h6C17: data_out = 8'h83;
                    16'h6C18: data_out = 8'h84;
                    16'h6C19: data_out = 8'h85;
                    16'h6C1A: data_out = 8'h86;
                    16'h6C1B: data_out = 8'h87;
                    16'h6C1C: data_out = 8'h88;
                    16'h6C1D: data_out = 8'h89;
                    16'h6C1E: data_out = 8'h8A;
                    16'h6C1F: data_out = 8'h8B;
                    16'h6C20: data_out = 8'h8C;
                    16'h6C21: data_out = 8'h8D;
                    16'h6C22: data_out = 8'h8E;
                    16'h6C23: data_out = 8'h8F;
                    16'h6C24: data_out = 8'h90;
                    16'h6C25: data_out = 8'h91;
                    16'h6C26: data_out = 8'h92;
                    16'h6C27: data_out = 8'h93;
                    16'h6C28: data_out = 8'h94;
                    16'h6C29: data_out = 8'h95;
                    16'h6C2A: data_out = 8'h96;
                    16'h6C2B: data_out = 8'h97;
                    16'h6C2C: data_out = 8'h98;
                    16'h6C2D: data_out = 8'h99;
                    16'h6C2E: data_out = 8'h9A;
                    16'h6C2F: data_out = 8'h9B;
                    16'h6C30: data_out = 8'h9C;
                    16'h6C31: data_out = 8'h9D;
                    16'h6C32: data_out = 8'h9E;
                    16'h6C33: data_out = 8'h9F;
                    16'h6C34: data_out = 8'hA0;
                    16'h6C35: data_out = 8'hA1;
                    16'h6C36: data_out = 8'hA2;
                    16'h6C37: data_out = 8'hA3;
                    16'h6C38: data_out = 8'hA4;
                    16'h6C39: data_out = 8'hA5;
                    16'h6C3A: data_out = 8'hA6;
                    16'h6C3B: data_out = 8'hA7;
                    16'h6C3C: data_out = 8'hA8;
                    16'h6C3D: data_out = 8'hA9;
                    16'h6C3E: data_out = 8'hAA;
                    16'h6C3F: data_out = 8'hAB;
                    16'h6C40: data_out = 8'hAC;
                    16'h6C41: data_out = 8'hAD;
                    16'h6C42: data_out = 8'hAE;
                    16'h6C43: data_out = 8'hAF;
                    16'h6C44: data_out = 8'hB0;
                    16'h6C45: data_out = 8'hB1;
                    16'h6C46: data_out = 8'hB2;
                    16'h6C47: data_out = 8'hB3;
                    16'h6C48: data_out = 8'hB4;
                    16'h6C49: data_out = 8'hB5;
                    16'h6C4A: data_out = 8'hB6;
                    16'h6C4B: data_out = 8'hB7;
                    16'h6C4C: data_out = 8'hB8;
                    16'h6C4D: data_out = 8'hB9;
                    16'h6C4E: data_out = 8'hBA;
                    16'h6C4F: data_out = 8'hBB;
                    16'h6C50: data_out = 8'hBC;
                    16'h6C51: data_out = 8'hBD;
                    16'h6C52: data_out = 8'hBE;
                    16'h6C53: data_out = 8'hBF;
                    16'h6C54: data_out = 8'hC0;
                    16'h6C55: data_out = 8'hC1;
                    16'h6C56: data_out = 8'hC2;
                    16'h6C57: data_out = 8'hC3;
                    16'h6C58: data_out = 8'hC4;
                    16'h6C59: data_out = 8'hC5;
                    16'h6C5A: data_out = 8'hC6;
                    16'h6C5B: data_out = 8'hC7;
                    16'h6C5C: data_out = 8'hC8;
                    16'h6C5D: data_out = 8'hC9;
                    16'h6C5E: data_out = 8'hCA;
                    16'h6C5F: data_out = 8'hCB;
                    16'h6C60: data_out = 8'hCC;
                    16'h6C61: data_out = 8'hCD;
                    16'h6C62: data_out = 8'hCE;
                    16'h6C63: data_out = 8'hCF;
                    16'h6C64: data_out = 8'hD0;
                    16'h6C65: data_out = 8'hD1;
                    16'h6C66: data_out = 8'hD2;
                    16'h6C67: data_out = 8'hD3;
                    16'h6C68: data_out = 8'hD4;
                    16'h6C69: data_out = 8'hD5;
                    16'h6C6A: data_out = 8'hD6;
                    16'h6C6B: data_out = 8'hD7;
                    16'h6C6C: data_out = 8'hD8;
                    16'h6C6D: data_out = 8'hD9;
                    16'h6C6E: data_out = 8'hDA;
                    16'h6C6F: data_out = 8'hDB;
                    16'h6C70: data_out = 8'hDC;
                    16'h6C71: data_out = 8'hDD;
                    16'h6C72: data_out = 8'hDE;
                    16'h6C73: data_out = 8'hDF;
                    16'h6C74: data_out = 8'hE0;
                    16'h6C75: data_out = 8'hE1;
                    16'h6C76: data_out = 8'hE2;
                    16'h6C77: data_out = 8'hE3;
                    16'h6C78: data_out = 8'hE4;
                    16'h6C79: data_out = 8'hE5;
                    16'h6C7A: data_out = 8'hE6;
                    16'h6C7B: data_out = 8'hE7;
                    16'h6C7C: data_out = 8'hE8;
                    16'h6C7D: data_out = 8'hE9;
                    16'h6C7E: data_out = 8'hEA;
                    16'h6C7F: data_out = 8'hEB;
                    16'h6C80: data_out = 8'h6C;
                    16'h6C81: data_out = 8'h6B;
                    16'h6C82: data_out = 8'h6A;
                    16'h6C83: data_out = 8'h69;
                    16'h6C84: data_out = 8'h68;
                    16'h6C85: data_out = 8'h67;
                    16'h6C86: data_out = 8'h66;
                    16'h6C87: data_out = 8'h65;
                    16'h6C88: data_out = 8'h64;
                    16'h6C89: data_out = 8'h63;
                    16'h6C8A: data_out = 8'h62;
                    16'h6C8B: data_out = 8'h61;
                    16'h6C8C: data_out = 8'h60;
                    16'h6C8D: data_out = 8'h5F;
                    16'h6C8E: data_out = 8'h5E;
                    16'h6C8F: data_out = 8'h5D;
                    16'h6C90: data_out = 8'h5C;
                    16'h6C91: data_out = 8'h5B;
                    16'h6C92: data_out = 8'h5A;
                    16'h6C93: data_out = 8'h59;
                    16'h6C94: data_out = 8'h58;
                    16'h6C95: data_out = 8'h57;
                    16'h6C96: data_out = 8'h56;
                    16'h6C97: data_out = 8'h55;
                    16'h6C98: data_out = 8'h54;
                    16'h6C99: data_out = 8'h53;
                    16'h6C9A: data_out = 8'h52;
                    16'h6C9B: data_out = 8'h51;
                    16'h6C9C: data_out = 8'h50;
                    16'h6C9D: data_out = 8'h4F;
                    16'h6C9E: data_out = 8'h4E;
                    16'h6C9F: data_out = 8'h4D;
                    16'h6CA0: data_out = 8'h4C;
                    16'h6CA1: data_out = 8'h4B;
                    16'h6CA2: data_out = 8'h4A;
                    16'h6CA3: data_out = 8'h49;
                    16'h6CA4: data_out = 8'h48;
                    16'h6CA5: data_out = 8'h47;
                    16'h6CA6: data_out = 8'h46;
                    16'h6CA7: data_out = 8'h45;
                    16'h6CA8: data_out = 8'h44;
                    16'h6CA9: data_out = 8'h43;
                    16'h6CAA: data_out = 8'h42;
                    16'h6CAB: data_out = 8'h41;
                    16'h6CAC: data_out = 8'h40;
                    16'h6CAD: data_out = 8'h3F;
                    16'h6CAE: data_out = 8'h3E;
                    16'h6CAF: data_out = 8'h3D;
                    16'h6CB0: data_out = 8'h3C;
                    16'h6CB1: data_out = 8'h3B;
                    16'h6CB2: data_out = 8'h3A;
                    16'h6CB3: data_out = 8'h39;
                    16'h6CB4: data_out = 8'h38;
                    16'h6CB5: data_out = 8'h37;
                    16'h6CB6: data_out = 8'h36;
                    16'h6CB7: data_out = 8'h35;
                    16'h6CB8: data_out = 8'h34;
                    16'h6CB9: data_out = 8'h33;
                    16'h6CBA: data_out = 8'h32;
                    16'h6CBB: data_out = 8'h31;
                    16'h6CBC: data_out = 8'h30;
                    16'h6CBD: data_out = 8'h2F;
                    16'h6CBE: data_out = 8'h2E;
                    16'h6CBF: data_out = 8'h2D;
                    16'h6CC0: data_out = 8'h2C;
                    16'h6CC1: data_out = 8'h2B;
                    16'h6CC2: data_out = 8'h2A;
                    16'h6CC3: data_out = 8'h29;
                    16'h6CC4: data_out = 8'h28;
                    16'h6CC5: data_out = 8'h27;
                    16'h6CC6: data_out = 8'h26;
                    16'h6CC7: data_out = 8'h25;
                    16'h6CC8: data_out = 8'h24;
                    16'h6CC9: data_out = 8'h23;
                    16'h6CCA: data_out = 8'h22;
                    16'h6CCB: data_out = 8'h21;
                    16'h6CCC: data_out = 8'h20;
                    16'h6CCD: data_out = 8'h1F;
                    16'h6CCE: data_out = 8'h1E;
                    16'h6CCF: data_out = 8'h1D;
                    16'h6CD0: data_out = 8'h1C;
                    16'h6CD1: data_out = 8'h1B;
                    16'h6CD2: data_out = 8'h1A;
                    16'h6CD3: data_out = 8'h19;
                    16'h6CD4: data_out = 8'h18;
                    16'h6CD5: data_out = 8'h17;
                    16'h6CD6: data_out = 8'h16;
                    16'h6CD7: data_out = 8'h15;
                    16'h6CD8: data_out = 8'h14;
                    16'h6CD9: data_out = 8'h13;
                    16'h6CDA: data_out = 8'h12;
                    16'h6CDB: data_out = 8'h11;
                    16'h6CDC: data_out = 8'h10;
                    16'h6CDD: data_out = 8'hF;
                    16'h6CDE: data_out = 8'hE;
                    16'h6CDF: data_out = 8'hD;
                    16'h6CE0: data_out = 8'hC;
                    16'h6CE1: data_out = 8'hB;
                    16'h6CE2: data_out = 8'hA;
                    16'h6CE3: data_out = 8'h9;
                    16'h6CE4: data_out = 8'h8;
                    16'h6CE5: data_out = 8'h7;
                    16'h6CE6: data_out = 8'h6;
                    16'h6CE7: data_out = 8'h5;
                    16'h6CE8: data_out = 8'h4;
                    16'h6CE9: data_out = 8'h3;
                    16'h6CEA: data_out = 8'h2;
                    16'h6CEB: data_out = 8'h1;
                    16'h6CEC: data_out = 8'h0;
                    16'h6CED: data_out = 8'h81;
                    16'h6CEE: data_out = 8'h82;
                    16'h6CEF: data_out = 8'h83;
                    16'h6CF0: data_out = 8'h84;
                    16'h6CF1: data_out = 8'h85;
                    16'h6CF2: data_out = 8'h86;
                    16'h6CF3: data_out = 8'h87;
                    16'h6CF4: data_out = 8'h88;
                    16'h6CF5: data_out = 8'h89;
                    16'h6CF6: data_out = 8'h8A;
                    16'h6CF7: data_out = 8'h8B;
                    16'h6CF8: data_out = 8'h8C;
                    16'h6CF9: data_out = 8'h8D;
                    16'h6CFA: data_out = 8'h8E;
                    16'h6CFB: data_out = 8'h8F;
                    16'h6CFC: data_out = 8'h90;
                    16'h6CFD: data_out = 8'h91;
                    16'h6CFE: data_out = 8'h92;
                    16'h6CFF: data_out = 8'h93;
                    16'h6D00: data_out = 8'h6D;
                    16'h6D01: data_out = 8'h6E;
                    16'h6D02: data_out = 8'h6F;
                    16'h6D03: data_out = 8'h70;
                    16'h6D04: data_out = 8'h71;
                    16'h6D05: data_out = 8'h72;
                    16'h6D06: data_out = 8'h73;
                    16'h6D07: data_out = 8'h74;
                    16'h6D08: data_out = 8'h75;
                    16'h6D09: data_out = 8'h76;
                    16'h6D0A: data_out = 8'h77;
                    16'h6D0B: data_out = 8'h78;
                    16'h6D0C: data_out = 8'h79;
                    16'h6D0D: data_out = 8'h7A;
                    16'h6D0E: data_out = 8'h7B;
                    16'h6D0F: data_out = 8'h7C;
                    16'h6D10: data_out = 8'h7D;
                    16'h6D11: data_out = 8'h7E;
                    16'h6D12: data_out = 8'h7F;
                    16'h6D13: data_out = 8'h80;
                    16'h6D14: data_out = 8'h81;
                    16'h6D15: data_out = 8'h82;
                    16'h6D16: data_out = 8'h83;
                    16'h6D17: data_out = 8'h84;
                    16'h6D18: data_out = 8'h85;
                    16'h6D19: data_out = 8'h86;
                    16'h6D1A: data_out = 8'h87;
                    16'h6D1B: data_out = 8'h88;
                    16'h6D1C: data_out = 8'h89;
                    16'h6D1D: data_out = 8'h8A;
                    16'h6D1E: data_out = 8'h8B;
                    16'h6D1F: data_out = 8'h8C;
                    16'h6D20: data_out = 8'h8D;
                    16'h6D21: data_out = 8'h8E;
                    16'h6D22: data_out = 8'h8F;
                    16'h6D23: data_out = 8'h90;
                    16'h6D24: data_out = 8'h91;
                    16'h6D25: data_out = 8'h92;
                    16'h6D26: data_out = 8'h93;
                    16'h6D27: data_out = 8'h94;
                    16'h6D28: data_out = 8'h95;
                    16'h6D29: data_out = 8'h96;
                    16'h6D2A: data_out = 8'h97;
                    16'h6D2B: data_out = 8'h98;
                    16'h6D2C: data_out = 8'h99;
                    16'h6D2D: data_out = 8'h9A;
                    16'h6D2E: data_out = 8'h9B;
                    16'h6D2F: data_out = 8'h9C;
                    16'h6D30: data_out = 8'h9D;
                    16'h6D31: data_out = 8'h9E;
                    16'h6D32: data_out = 8'h9F;
                    16'h6D33: data_out = 8'hA0;
                    16'h6D34: data_out = 8'hA1;
                    16'h6D35: data_out = 8'hA2;
                    16'h6D36: data_out = 8'hA3;
                    16'h6D37: data_out = 8'hA4;
                    16'h6D38: data_out = 8'hA5;
                    16'h6D39: data_out = 8'hA6;
                    16'h6D3A: data_out = 8'hA7;
                    16'h6D3B: data_out = 8'hA8;
                    16'h6D3C: data_out = 8'hA9;
                    16'h6D3D: data_out = 8'hAA;
                    16'h6D3E: data_out = 8'hAB;
                    16'h6D3F: data_out = 8'hAC;
                    16'h6D40: data_out = 8'hAD;
                    16'h6D41: data_out = 8'hAE;
                    16'h6D42: data_out = 8'hAF;
                    16'h6D43: data_out = 8'hB0;
                    16'h6D44: data_out = 8'hB1;
                    16'h6D45: data_out = 8'hB2;
                    16'h6D46: data_out = 8'hB3;
                    16'h6D47: data_out = 8'hB4;
                    16'h6D48: data_out = 8'hB5;
                    16'h6D49: data_out = 8'hB6;
                    16'h6D4A: data_out = 8'hB7;
                    16'h6D4B: data_out = 8'hB8;
                    16'h6D4C: data_out = 8'hB9;
                    16'h6D4D: data_out = 8'hBA;
                    16'h6D4E: data_out = 8'hBB;
                    16'h6D4F: data_out = 8'hBC;
                    16'h6D50: data_out = 8'hBD;
                    16'h6D51: data_out = 8'hBE;
                    16'h6D52: data_out = 8'hBF;
                    16'h6D53: data_out = 8'hC0;
                    16'h6D54: data_out = 8'hC1;
                    16'h6D55: data_out = 8'hC2;
                    16'h6D56: data_out = 8'hC3;
                    16'h6D57: data_out = 8'hC4;
                    16'h6D58: data_out = 8'hC5;
                    16'h6D59: data_out = 8'hC6;
                    16'h6D5A: data_out = 8'hC7;
                    16'h6D5B: data_out = 8'hC8;
                    16'h6D5C: data_out = 8'hC9;
                    16'h6D5D: data_out = 8'hCA;
                    16'h6D5E: data_out = 8'hCB;
                    16'h6D5F: data_out = 8'hCC;
                    16'h6D60: data_out = 8'hCD;
                    16'h6D61: data_out = 8'hCE;
                    16'h6D62: data_out = 8'hCF;
                    16'h6D63: data_out = 8'hD0;
                    16'h6D64: data_out = 8'hD1;
                    16'h6D65: data_out = 8'hD2;
                    16'h6D66: data_out = 8'hD3;
                    16'h6D67: data_out = 8'hD4;
                    16'h6D68: data_out = 8'hD5;
                    16'h6D69: data_out = 8'hD6;
                    16'h6D6A: data_out = 8'hD7;
                    16'h6D6B: data_out = 8'hD8;
                    16'h6D6C: data_out = 8'hD9;
                    16'h6D6D: data_out = 8'hDA;
                    16'h6D6E: data_out = 8'hDB;
                    16'h6D6F: data_out = 8'hDC;
                    16'h6D70: data_out = 8'hDD;
                    16'h6D71: data_out = 8'hDE;
                    16'h6D72: data_out = 8'hDF;
                    16'h6D73: data_out = 8'hE0;
                    16'h6D74: data_out = 8'hE1;
                    16'h6D75: data_out = 8'hE2;
                    16'h6D76: data_out = 8'hE3;
                    16'h6D77: data_out = 8'hE4;
                    16'h6D78: data_out = 8'hE5;
                    16'h6D79: data_out = 8'hE6;
                    16'h6D7A: data_out = 8'hE7;
                    16'h6D7B: data_out = 8'hE8;
                    16'h6D7C: data_out = 8'hE9;
                    16'h6D7D: data_out = 8'hEA;
                    16'h6D7E: data_out = 8'hEB;
                    16'h6D7F: data_out = 8'hEC;
                    16'h6D80: data_out = 8'h6D;
                    16'h6D81: data_out = 8'h6C;
                    16'h6D82: data_out = 8'h6B;
                    16'h6D83: data_out = 8'h6A;
                    16'h6D84: data_out = 8'h69;
                    16'h6D85: data_out = 8'h68;
                    16'h6D86: data_out = 8'h67;
                    16'h6D87: data_out = 8'h66;
                    16'h6D88: data_out = 8'h65;
                    16'h6D89: data_out = 8'h64;
                    16'h6D8A: data_out = 8'h63;
                    16'h6D8B: data_out = 8'h62;
                    16'h6D8C: data_out = 8'h61;
                    16'h6D8D: data_out = 8'h60;
                    16'h6D8E: data_out = 8'h5F;
                    16'h6D8F: data_out = 8'h5E;
                    16'h6D90: data_out = 8'h5D;
                    16'h6D91: data_out = 8'h5C;
                    16'h6D92: data_out = 8'h5B;
                    16'h6D93: data_out = 8'h5A;
                    16'h6D94: data_out = 8'h59;
                    16'h6D95: data_out = 8'h58;
                    16'h6D96: data_out = 8'h57;
                    16'h6D97: data_out = 8'h56;
                    16'h6D98: data_out = 8'h55;
                    16'h6D99: data_out = 8'h54;
                    16'h6D9A: data_out = 8'h53;
                    16'h6D9B: data_out = 8'h52;
                    16'h6D9C: data_out = 8'h51;
                    16'h6D9D: data_out = 8'h50;
                    16'h6D9E: data_out = 8'h4F;
                    16'h6D9F: data_out = 8'h4E;
                    16'h6DA0: data_out = 8'h4D;
                    16'h6DA1: data_out = 8'h4C;
                    16'h6DA2: data_out = 8'h4B;
                    16'h6DA3: data_out = 8'h4A;
                    16'h6DA4: data_out = 8'h49;
                    16'h6DA5: data_out = 8'h48;
                    16'h6DA6: data_out = 8'h47;
                    16'h6DA7: data_out = 8'h46;
                    16'h6DA8: data_out = 8'h45;
                    16'h6DA9: data_out = 8'h44;
                    16'h6DAA: data_out = 8'h43;
                    16'h6DAB: data_out = 8'h42;
                    16'h6DAC: data_out = 8'h41;
                    16'h6DAD: data_out = 8'h40;
                    16'h6DAE: data_out = 8'h3F;
                    16'h6DAF: data_out = 8'h3E;
                    16'h6DB0: data_out = 8'h3D;
                    16'h6DB1: data_out = 8'h3C;
                    16'h6DB2: data_out = 8'h3B;
                    16'h6DB3: data_out = 8'h3A;
                    16'h6DB4: data_out = 8'h39;
                    16'h6DB5: data_out = 8'h38;
                    16'h6DB6: data_out = 8'h37;
                    16'h6DB7: data_out = 8'h36;
                    16'h6DB8: data_out = 8'h35;
                    16'h6DB9: data_out = 8'h34;
                    16'h6DBA: data_out = 8'h33;
                    16'h6DBB: data_out = 8'h32;
                    16'h6DBC: data_out = 8'h31;
                    16'h6DBD: data_out = 8'h30;
                    16'h6DBE: data_out = 8'h2F;
                    16'h6DBF: data_out = 8'h2E;
                    16'h6DC0: data_out = 8'h2D;
                    16'h6DC1: data_out = 8'h2C;
                    16'h6DC2: data_out = 8'h2B;
                    16'h6DC3: data_out = 8'h2A;
                    16'h6DC4: data_out = 8'h29;
                    16'h6DC5: data_out = 8'h28;
                    16'h6DC6: data_out = 8'h27;
                    16'h6DC7: data_out = 8'h26;
                    16'h6DC8: data_out = 8'h25;
                    16'h6DC9: data_out = 8'h24;
                    16'h6DCA: data_out = 8'h23;
                    16'h6DCB: data_out = 8'h22;
                    16'h6DCC: data_out = 8'h21;
                    16'h6DCD: data_out = 8'h20;
                    16'h6DCE: data_out = 8'h1F;
                    16'h6DCF: data_out = 8'h1E;
                    16'h6DD0: data_out = 8'h1D;
                    16'h6DD1: data_out = 8'h1C;
                    16'h6DD2: data_out = 8'h1B;
                    16'h6DD3: data_out = 8'h1A;
                    16'h6DD4: data_out = 8'h19;
                    16'h6DD5: data_out = 8'h18;
                    16'h6DD6: data_out = 8'h17;
                    16'h6DD7: data_out = 8'h16;
                    16'h6DD8: data_out = 8'h15;
                    16'h6DD9: data_out = 8'h14;
                    16'h6DDA: data_out = 8'h13;
                    16'h6DDB: data_out = 8'h12;
                    16'h6DDC: data_out = 8'h11;
                    16'h6DDD: data_out = 8'h10;
                    16'h6DDE: data_out = 8'hF;
                    16'h6DDF: data_out = 8'hE;
                    16'h6DE0: data_out = 8'hD;
                    16'h6DE1: data_out = 8'hC;
                    16'h6DE2: data_out = 8'hB;
                    16'h6DE3: data_out = 8'hA;
                    16'h6DE4: data_out = 8'h9;
                    16'h6DE5: data_out = 8'h8;
                    16'h6DE6: data_out = 8'h7;
                    16'h6DE7: data_out = 8'h6;
                    16'h6DE8: data_out = 8'h5;
                    16'h6DE9: data_out = 8'h4;
                    16'h6DEA: data_out = 8'h3;
                    16'h6DEB: data_out = 8'h2;
                    16'h6DEC: data_out = 8'h1;
                    16'h6DED: data_out = 8'h0;
                    16'h6DEE: data_out = 8'h81;
                    16'h6DEF: data_out = 8'h82;
                    16'h6DF0: data_out = 8'h83;
                    16'h6DF1: data_out = 8'h84;
                    16'h6DF2: data_out = 8'h85;
                    16'h6DF3: data_out = 8'h86;
                    16'h6DF4: data_out = 8'h87;
                    16'h6DF5: data_out = 8'h88;
                    16'h6DF6: data_out = 8'h89;
                    16'h6DF7: data_out = 8'h8A;
                    16'h6DF8: data_out = 8'h8B;
                    16'h6DF9: data_out = 8'h8C;
                    16'h6DFA: data_out = 8'h8D;
                    16'h6DFB: data_out = 8'h8E;
                    16'h6DFC: data_out = 8'h8F;
                    16'h6DFD: data_out = 8'h90;
                    16'h6DFE: data_out = 8'h91;
                    16'h6DFF: data_out = 8'h92;
                    16'h6E00: data_out = 8'h6E;
                    16'h6E01: data_out = 8'h6F;
                    16'h6E02: data_out = 8'h70;
                    16'h6E03: data_out = 8'h71;
                    16'h6E04: data_out = 8'h72;
                    16'h6E05: data_out = 8'h73;
                    16'h6E06: data_out = 8'h74;
                    16'h6E07: data_out = 8'h75;
                    16'h6E08: data_out = 8'h76;
                    16'h6E09: data_out = 8'h77;
                    16'h6E0A: data_out = 8'h78;
                    16'h6E0B: data_out = 8'h79;
                    16'h6E0C: data_out = 8'h7A;
                    16'h6E0D: data_out = 8'h7B;
                    16'h6E0E: data_out = 8'h7C;
                    16'h6E0F: data_out = 8'h7D;
                    16'h6E10: data_out = 8'h7E;
                    16'h6E11: data_out = 8'h7F;
                    16'h6E12: data_out = 8'h80;
                    16'h6E13: data_out = 8'h81;
                    16'h6E14: data_out = 8'h82;
                    16'h6E15: data_out = 8'h83;
                    16'h6E16: data_out = 8'h84;
                    16'h6E17: data_out = 8'h85;
                    16'h6E18: data_out = 8'h86;
                    16'h6E19: data_out = 8'h87;
                    16'h6E1A: data_out = 8'h88;
                    16'h6E1B: data_out = 8'h89;
                    16'h6E1C: data_out = 8'h8A;
                    16'h6E1D: data_out = 8'h8B;
                    16'h6E1E: data_out = 8'h8C;
                    16'h6E1F: data_out = 8'h8D;
                    16'h6E20: data_out = 8'h8E;
                    16'h6E21: data_out = 8'h8F;
                    16'h6E22: data_out = 8'h90;
                    16'h6E23: data_out = 8'h91;
                    16'h6E24: data_out = 8'h92;
                    16'h6E25: data_out = 8'h93;
                    16'h6E26: data_out = 8'h94;
                    16'h6E27: data_out = 8'h95;
                    16'h6E28: data_out = 8'h96;
                    16'h6E29: data_out = 8'h97;
                    16'h6E2A: data_out = 8'h98;
                    16'h6E2B: data_out = 8'h99;
                    16'h6E2C: data_out = 8'h9A;
                    16'h6E2D: data_out = 8'h9B;
                    16'h6E2E: data_out = 8'h9C;
                    16'h6E2F: data_out = 8'h9D;
                    16'h6E30: data_out = 8'h9E;
                    16'h6E31: data_out = 8'h9F;
                    16'h6E32: data_out = 8'hA0;
                    16'h6E33: data_out = 8'hA1;
                    16'h6E34: data_out = 8'hA2;
                    16'h6E35: data_out = 8'hA3;
                    16'h6E36: data_out = 8'hA4;
                    16'h6E37: data_out = 8'hA5;
                    16'h6E38: data_out = 8'hA6;
                    16'h6E39: data_out = 8'hA7;
                    16'h6E3A: data_out = 8'hA8;
                    16'h6E3B: data_out = 8'hA9;
                    16'h6E3C: data_out = 8'hAA;
                    16'h6E3D: data_out = 8'hAB;
                    16'h6E3E: data_out = 8'hAC;
                    16'h6E3F: data_out = 8'hAD;
                    16'h6E40: data_out = 8'hAE;
                    16'h6E41: data_out = 8'hAF;
                    16'h6E42: data_out = 8'hB0;
                    16'h6E43: data_out = 8'hB1;
                    16'h6E44: data_out = 8'hB2;
                    16'h6E45: data_out = 8'hB3;
                    16'h6E46: data_out = 8'hB4;
                    16'h6E47: data_out = 8'hB5;
                    16'h6E48: data_out = 8'hB6;
                    16'h6E49: data_out = 8'hB7;
                    16'h6E4A: data_out = 8'hB8;
                    16'h6E4B: data_out = 8'hB9;
                    16'h6E4C: data_out = 8'hBA;
                    16'h6E4D: data_out = 8'hBB;
                    16'h6E4E: data_out = 8'hBC;
                    16'h6E4F: data_out = 8'hBD;
                    16'h6E50: data_out = 8'hBE;
                    16'h6E51: data_out = 8'hBF;
                    16'h6E52: data_out = 8'hC0;
                    16'h6E53: data_out = 8'hC1;
                    16'h6E54: data_out = 8'hC2;
                    16'h6E55: data_out = 8'hC3;
                    16'h6E56: data_out = 8'hC4;
                    16'h6E57: data_out = 8'hC5;
                    16'h6E58: data_out = 8'hC6;
                    16'h6E59: data_out = 8'hC7;
                    16'h6E5A: data_out = 8'hC8;
                    16'h6E5B: data_out = 8'hC9;
                    16'h6E5C: data_out = 8'hCA;
                    16'h6E5D: data_out = 8'hCB;
                    16'h6E5E: data_out = 8'hCC;
                    16'h6E5F: data_out = 8'hCD;
                    16'h6E60: data_out = 8'hCE;
                    16'h6E61: data_out = 8'hCF;
                    16'h6E62: data_out = 8'hD0;
                    16'h6E63: data_out = 8'hD1;
                    16'h6E64: data_out = 8'hD2;
                    16'h6E65: data_out = 8'hD3;
                    16'h6E66: data_out = 8'hD4;
                    16'h6E67: data_out = 8'hD5;
                    16'h6E68: data_out = 8'hD6;
                    16'h6E69: data_out = 8'hD7;
                    16'h6E6A: data_out = 8'hD8;
                    16'h6E6B: data_out = 8'hD9;
                    16'h6E6C: data_out = 8'hDA;
                    16'h6E6D: data_out = 8'hDB;
                    16'h6E6E: data_out = 8'hDC;
                    16'h6E6F: data_out = 8'hDD;
                    16'h6E70: data_out = 8'hDE;
                    16'h6E71: data_out = 8'hDF;
                    16'h6E72: data_out = 8'hE0;
                    16'h6E73: data_out = 8'hE1;
                    16'h6E74: data_out = 8'hE2;
                    16'h6E75: data_out = 8'hE3;
                    16'h6E76: data_out = 8'hE4;
                    16'h6E77: data_out = 8'hE5;
                    16'h6E78: data_out = 8'hE6;
                    16'h6E79: data_out = 8'hE7;
                    16'h6E7A: data_out = 8'hE8;
                    16'h6E7B: data_out = 8'hE9;
                    16'h6E7C: data_out = 8'hEA;
                    16'h6E7D: data_out = 8'hEB;
                    16'h6E7E: data_out = 8'hEC;
                    16'h6E7F: data_out = 8'hED;
                    16'h6E80: data_out = 8'h6E;
                    16'h6E81: data_out = 8'h6D;
                    16'h6E82: data_out = 8'h6C;
                    16'h6E83: data_out = 8'h6B;
                    16'h6E84: data_out = 8'h6A;
                    16'h6E85: data_out = 8'h69;
                    16'h6E86: data_out = 8'h68;
                    16'h6E87: data_out = 8'h67;
                    16'h6E88: data_out = 8'h66;
                    16'h6E89: data_out = 8'h65;
                    16'h6E8A: data_out = 8'h64;
                    16'h6E8B: data_out = 8'h63;
                    16'h6E8C: data_out = 8'h62;
                    16'h6E8D: data_out = 8'h61;
                    16'h6E8E: data_out = 8'h60;
                    16'h6E8F: data_out = 8'h5F;
                    16'h6E90: data_out = 8'h5E;
                    16'h6E91: data_out = 8'h5D;
                    16'h6E92: data_out = 8'h5C;
                    16'h6E93: data_out = 8'h5B;
                    16'h6E94: data_out = 8'h5A;
                    16'h6E95: data_out = 8'h59;
                    16'h6E96: data_out = 8'h58;
                    16'h6E97: data_out = 8'h57;
                    16'h6E98: data_out = 8'h56;
                    16'h6E99: data_out = 8'h55;
                    16'h6E9A: data_out = 8'h54;
                    16'h6E9B: data_out = 8'h53;
                    16'h6E9C: data_out = 8'h52;
                    16'h6E9D: data_out = 8'h51;
                    16'h6E9E: data_out = 8'h50;
                    16'h6E9F: data_out = 8'h4F;
                    16'h6EA0: data_out = 8'h4E;
                    16'h6EA1: data_out = 8'h4D;
                    16'h6EA2: data_out = 8'h4C;
                    16'h6EA3: data_out = 8'h4B;
                    16'h6EA4: data_out = 8'h4A;
                    16'h6EA5: data_out = 8'h49;
                    16'h6EA6: data_out = 8'h48;
                    16'h6EA7: data_out = 8'h47;
                    16'h6EA8: data_out = 8'h46;
                    16'h6EA9: data_out = 8'h45;
                    16'h6EAA: data_out = 8'h44;
                    16'h6EAB: data_out = 8'h43;
                    16'h6EAC: data_out = 8'h42;
                    16'h6EAD: data_out = 8'h41;
                    16'h6EAE: data_out = 8'h40;
                    16'h6EAF: data_out = 8'h3F;
                    16'h6EB0: data_out = 8'h3E;
                    16'h6EB1: data_out = 8'h3D;
                    16'h6EB2: data_out = 8'h3C;
                    16'h6EB3: data_out = 8'h3B;
                    16'h6EB4: data_out = 8'h3A;
                    16'h6EB5: data_out = 8'h39;
                    16'h6EB6: data_out = 8'h38;
                    16'h6EB7: data_out = 8'h37;
                    16'h6EB8: data_out = 8'h36;
                    16'h6EB9: data_out = 8'h35;
                    16'h6EBA: data_out = 8'h34;
                    16'h6EBB: data_out = 8'h33;
                    16'h6EBC: data_out = 8'h32;
                    16'h6EBD: data_out = 8'h31;
                    16'h6EBE: data_out = 8'h30;
                    16'h6EBF: data_out = 8'h2F;
                    16'h6EC0: data_out = 8'h2E;
                    16'h6EC1: data_out = 8'h2D;
                    16'h6EC2: data_out = 8'h2C;
                    16'h6EC3: data_out = 8'h2B;
                    16'h6EC4: data_out = 8'h2A;
                    16'h6EC5: data_out = 8'h29;
                    16'h6EC6: data_out = 8'h28;
                    16'h6EC7: data_out = 8'h27;
                    16'h6EC8: data_out = 8'h26;
                    16'h6EC9: data_out = 8'h25;
                    16'h6ECA: data_out = 8'h24;
                    16'h6ECB: data_out = 8'h23;
                    16'h6ECC: data_out = 8'h22;
                    16'h6ECD: data_out = 8'h21;
                    16'h6ECE: data_out = 8'h20;
                    16'h6ECF: data_out = 8'h1F;
                    16'h6ED0: data_out = 8'h1E;
                    16'h6ED1: data_out = 8'h1D;
                    16'h6ED2: data_out = 8'h1C;
                    16'h6ED3: data_out = 8'h1B;
                    16'h6ED4: data_out = 8'h1A;
                    16'h6ED5: data_out = 8'h19;
                    16'h6ED6: data_out = 8'h18;
                    16'h6ED7: data_out = 8'h17;
                    16'h6ED8: data_out = 8'h16;
                    16'h6ED9: data_out = 8'h15;
                    16'h6EDA: data_out = 8'h14;
                    16'h6EDB: data_out = 8'h13;
                    16'h6EDC: data_out = 8'h12;
                    16'h6EDD: data_out = 8'h11;
                    16'h6EDE: data_out = 8'h10;
                    16'h6EDF: data_out = 8'hF;
                    16'h6EE0: data_out = 8'hE;
                    16'h6EE1: data_out = 8'hD;
                    16'h6EE2: data_out = 8'hC;
                    16'h6EE3: data_out = 8'hB;
                    16'h6EE4: data_out = 8'hA;
                    16'h6EE5: data_out = 8'h9;
                    16'h6EE6: data_out = 8'h8;
                    16'h6EE7: data_out = 8'h7;
                    16'h6EE8: data_out = 8'h6;
                    16'h6EE9: data_out = 8'h5;
                    16'h6EEA: data_out = 8'h4;
                    16'h6EEB: data_out = 8'h3;
                    16'h6EEC: data_out = 8'h2;
                    16'h6EED: data_out = 8'h1;
                    16'h6EEE: data_out = 8'h0;
                    16'h6EEF: data_out = 8'h81;
                    16'h6EF0: data_out = 8'h82;
                    16'h6EF1: data_out = 8'h83;
                    16'h6EF2: data_out = 8'h84;
                    16'h6EF3: data_out = 8'h85;
                    16'h6EF4: data_out = 8'h86;
                    16'h6EF5: data_out = 8'h87;
                    16'h6EF6: data_out = 8'h88;
                    16'h6EF7: data_out = 8'h89;
                    16'h6EF8: data_out = 8'h8A;
                    16'h6EF9: data_out = 8'h8B;
                    16'h6EFA: data_out = 8'h8C;
                    16'h6EFB: data_out = 8'h8D;
                    16'h6EFC: data_out = 8'h8E;
                    16'h6EFD: data_out = 8'h8F;
                    16'h6EFE: data_out = 8'h90;
                    16'h6EFF: data_out = 8'h91;
                    16'h6F00: data_out = 8'h6F;
                    16'h6F01: data_out = 8'h70;
                    16'h6F02: data_out = 8'h71;
                    16'h6F03: data_out = 8'h72;
                    16'h6F04: data_out = 8'h73;
                    16'h6F05: data_out = 8'h74;
                    16'h6F06: data_out = 8'h75;
                    16'h6F07: data_out = 8'h76;
                    16'h6F08: data_out = 8'h77;
                    16'h6F09: data_out = 8'h78;
                    16'h6F0A: data_out = 8'h79;
                    16'h6F0B: data_out = 8'h7A;
                    16'h6F0C: data_out = 8'h7B;
                    16'h6F0D: data_out = 8'h7C;
                    16'h6F0E: data_out = 8'h7D;
                    16'h6F0F: data_out = 8'h7E;
                    16'h6F10: data_out = 8'h7F;
                    16'h6F11: data_out = 8'h80;
                    16'h6F12: data_out = 8'h81;
                    16'h6F13: data_out = 8'h82;
                    16'h6F14: data_out = 8'h83;
                    16'h6F15: data_out = 8'h84;
                    16'h6F16: data_out = 8'h85;
                    16'h6F17: data_out = 8'h86;
                    16'h6F18: data_out = 8'h87;
                    16'h6F19: data_out = 8'h88;
                    16'h6F1A: data_out = 8'h89;
                    16'h6F1B: data_out = 8'h8A;
                    16'h6F1C: data_out = 8'h8B;
                    16'h6F1D: data_out = 8'h8C;
                    16'h6F1E: data_out = 8'h8D;
                    16'h6F1F: data_out = 8'h8E;
                    16'h6F20: data_out = 8'h8F;
                    16'h6F21: data_out = 8'h90;
                    16'h6F22: data_out = 8'h91;
                    16'h6F23: data_out = 8'h92;
                    16'h6F24: data_out = 8'h93;
                    16'h6F25: data_out = 8'h94;
                    16'h6F26: data_out = 8'h95;
                    16'h6F27: data_out = 8'h96;
                    16'h6F28: data_out = 8'h97;
                    16'h6F29: data_out = 8'h98;
                    16'h6F2A: data_out = 8'h99;
                    16'h6F2B: data_out = 8'h9A;
                    16'h6F2C: data_out = 8'h9B;
                    16'h6F2D: data_out = 8'h9C;
                    16'h6F2E: data_out = 8'h9D;
                    16'h6F2F: data_out = 8'h9E;
                    16'h6F30: data_out = 8'h9F;
                    16'h6F31: data_out = 8'hA0;
                    16'h6F32: data_out = 8'hA1;
                    16'h6F33: data_out = 8'hA2;
                    16'h6F34: data_out = 8'hA3;
                    16'h6F35: data_out = 8'hA4;
                    16'h6F36: data_out = 8'hA5;
                    16'h6F37: data_out = 8'hA6;
                    16'h6F38: data_out = 8'hA7;
                    16'h6F39: data_out = 8'hA8;
                    16'h6F3A: data_out = 8'hA9;
                    16'h6F3B: data_out = 8'hAA;
                    16'h6F3C: data_out = 8'hAB;
                    16'h6F3D: data_out = 8'hAC;
                    16'h6F3E: data_out = 8'hAD;
                    16'h6F3F: data_out = 8'hAE;
                    16'h6F40: data_out = 8'hAF;
                    16'h6F41: data_out = 8'hB0;
                    16'h6F42: data_out = 8'hB1;
                    16'h6F43: data_out = 8'hB2;
                    16'h6F44: data_out = 8'hB3;
                    16'h6F45: data_out = 8'hB4;
                    16'h6F46: data_out = 8'hB5;
                    16'h6F47: data_out = 8'hB6;
                    16'h6F48: data_out = 8'hB7;
                    16'h6F49: data_out = 8'hB8;
                    16'h6F4A: data_out = 8'hB9;
                    16'h6F4B: data_out = 8'hBA;
                    16'h6F4C: data_out = 8'hBB;
                    16'h6F4D: data_out = 8'hBC;
                    16'h6F4E: data_out = 8'hBD;
                    16'h6F4F: data_out = 8'hBE;
                    16'h6F50: data_out = 8'hBF;
                    16'h6F51: data_out = 8'hC0;
                    16'h6F52: data_out = 8'hC1;
                    16'h6F53: data_out = 8'hC2;
                    16'h6F54: data_out = 8'hC3;
                    16'h6F55: data_out = 8'hC4;
                    16'h6F56: data_out = 8'hC5;
                    16'h6F57: data_out = 8'hC6;
                    16'h6F58: data_out = 8'hC7;
                    16'h6F59: data_out = 8'hC8;
                    16'h6F5A: data_out = 8'hC9;
                    16'h6F5B: data_out = 8'hCA;
                    16'h6F5C: data_out = 8'hCB;
                    16'h6F5D: data_out = 8'hCC;
                    16'h6F5E: data_out = 8'hCD;
                    16'h6F5F: data_out = 8'hCE;
                    16'h6F60: data_out = 8'hCF;
                    16'h6F61: data_out = 8'hD0;
                    16'h6F62: data_out = 8'hD1;
                    16'h6F63: data_out = 8'hD2;
                    16'h6F64: data_out = 8'hD3;
                    16'h6F65: data_out = 8'hD4;
                    16'h6F66: data_out = 8'hD5;
                    16'h6F67: data_out = 8'hD6;
                    16'h6F68: data_out = 8'hD7;
                    16'h6F69: data_out = 8'hD8;
                    16'h6F6A: data_out = 8'hD9;
                    16'h6F6B: data_out = 8'hDA;
                    16'h6F6C: data_out = 8'hDB;
                    16'h6F6D: data_out = 8'hDC;
                    16'h6F6E: data_out = 8'hDD;
                    16'h6F6F: data_out = 8'hDE;
                    16'h6F70: data_out = 8'hDF;
                    16'h6F71: data_out = 8'hE0;
                    16'h6F72: data_out = 8'hE1;
                    16'h6F73: data_out = 8'hE2;
                    16'h6F74: data_out = 8'hE3;
                    16'h6F75: data_out = 8'hE4;
                    16'h6F76: data_out = 8'hE5;
                    16'h6F77: data_out = 8'hE6;
                    16'h6F78: data_out = 8'hE7;
                    16'h6F79: data_out = 8'hE8;
                    16'h6F7A: data_out = 8'hE9;
                    16'h6F7B: data_out = 8'hEA;
                    16'h6F7C: data_out = 8'hEB;
                    16'h6F7D: data_out = 8'hEC;
                    16'h6F7E: data_out = 8'hED;
                    16'h6F7F: data_out = 8'hEE;
                    16'h6F80: data_out = 8'h6F;
                    16'h6F81: data_out = 8'h6E;
                    16'h6F82: data_out = 8'h6D;
                    16'h6F83: data_out = 8'h6C;
                    16'h6F84: data_out = 8'h6B;
                    16'h6F85: data_out = 8'h6A;
                    16'h6F86: data_out = 8'h69;
                    16'h6F87: data_out = 8'h68;
                    16'h6F88: data_out = 8'h67;
                    16'h6F89: data_out = 8'h66;
                    16'h6F8A: data_out = 8'h65;
                    16'h6F8B: data_out = 8'h64;
                    16'h6F8C: data_out = 8'h63;
                    16'h6F8D: data_out = 8'h62;
                    16'h6F8E: data_out = 8'h61;
                    16'h6F8F: data_out = 8'h60;
                    16'h6F90: data_out = 8'h5F;
                    16'h6F91: data_out = 8'h5E;
                    16'h6F92: data_out = 8'h5D;
                    16'h6F93: data_out = 8'h5C;
                    16'h6F94: data_out = 8'h5B;
                    16'h6F95: data_out = 8'h5A;
                    16'h6F96: data_out = 8'h59;
                    16'h6F97: data_out = 8'h58;
                    16'h6F98: data_out = 8'h57;
                    16'h6F99: data_out = 8'h56;
                    16'h6F9A: data_out = 8'h55;
                    16'h6F9B: data_out = 8'h54;
                    16'h6F9C: data_out = 8'h53;
                    16'h6F9D: data_out = 8'h52;
                    16'h6F9E: data_out = 8'h51;
                    16'h6F9F: data_out = 8'h50;
                    16'h6FA0: data_out = 8'h4F;
                    16'h6FA1: data_out = 8'h4E;
                    16'h6FA2: data_out = 8'h4D;
                    16'h6FA3: data_out = 8'h4C;
                    16'h6FA4: data_out = 8'h4B;
                    16'h6FA5: data_out = 8'h4A;
                    16'h6FA6: data_out = 8'h49;
                    16'h6FA7: data_out = 8'h48;
                    16'h6FA8: data_out = 8'h47;
                    16'h6FA9: data_out = 8'h46;
                    16'h6FAA: data_out = 8'h45;
                    16'h6FAB: data_out = 8'h44;
                    16'h6FAC: data_out = 8'h43;
                    16'h6FAD: data_out = 8'h42;
                    16'h6FAE: data_out = 8'h41;
                    16'h6FAF: data_out = 8'h40;
                    16'h6FB0: data_out = 8'h3F;
                    16'h6FB1: data_out = 8'h3E;
                    16'h6FB2: data_out = 8'h3D;
                    16'h6FB3: data_out = 8'h3C;
                    16'h6FB4: data_out = 8'h3B;
                    16'h6FB5: data_out = 8'h3A;
                    16'h6FB6: data_out = 8'h39;
                    16'h6FB7: data_out = 8'h38;
                    16'h6FB8: data_out = 8'h37;
                    16'h6FB9: data_out = 8'h36;
                    16'h6FBA: data_out = 8'h35;
                    16'h6FBB: data_out = 8'h34;
                    16'h6FBC: data_out = 8'h33;
                    16'h6FBD: data_out = 8'h32;
                    16'h6FBE: data_out = 8'h31;
                    16'h6FBF: data_out = 8'h30;
                    16'h6FC0: data_out = 8'h2F;
                    16'h6FC1: data_out = 8'h2E;
                    16'h6FC2: data_out = 8'h2D;
                    16'h6FC3: data_out = 8'h2C;
                    16'h6FC4: data_out = 8'h2B;
                    16'h6FC5: data_out = 8'h2A;
                    16'h6FC6: data_out = 8'h29;
                    16'h6FC7: data_out = 8'h28;
                    16'h6FC8: data_out = 8'h27;
                    16'h6FC9: data_out = 8'h26;
                    16'h6FCA: data_out = 8'h25;
                    16'h6FCB: data_out = 8'h24;
                    16'h6FCC: data_out = 8'h23;
                    16'h6FCD: data_out = 8'h22;
                    16'h6FCE: data_out = 8'h21;
                    16'h6FCF: data_out = 8'h20;
                    16'h6FD0: data_out = 8'h1F;
                    16'h6FD1: data_out = 8'h1E;
                    16'h6FD2: data_out = 8'h1D;
                    16'h6FD3: data_out = 8'h1C;
                    16'h6FD4: data_out = 8'h1B;
                    16'h6FD5: data_out = 8'h1A;
                    16'h6FD6: data_out = 8'h19;
                    16'h6FD7: data_out = 8'h18;
                    16'h6FD8: data_out = 8'h17;
                    16'h6FD9: data_out = 8'h16;
                    16'h6FDA: data_out = 8'h15;
                    16'h6FDB: data_out = 8'h14;
                    16'h6FDC: data_out = 8'h13;
                    16'h6FDD: data_out = 8'h12;
                    16'h6FDE: data_out = 8'h11;
                    16'h6FDF: data_out = 8'h10;
                    16'h6FE0: data_out = 8'hF;
                    16'h6FE1: data_out = 8'hE;
                    16'h6FE2: data_out = 8'hD;
                    16'h6FE3: data_out = 8'hC;
                    16'h6FE4: data_out = 8'hB;
                    16'h6FE5: data_out = 8'hA;
                    16'h6FE6: data_out = 8'h9;
                    16'h6FE7: data_out = 8'h8;
                    16'h6FE8: data_out = 8'h7;
                    16'h6FE9: data_out = 8'h6;
                    16'h6FEA: data_out = 8'h5;
                    16'h6FEB: data_out = 8'h4;
                    16'h6FEC: data_out = 8'h3;
                    16'h6FED: data_out = 8'h2;
                    16'h6FEE: data_out = 8'h1;
                    16'h6FEF: data_out = 8'h0;
                    16'h6FF0: data_out = 8'h81;
                    16'h6FF1: data_out = 8'h82;
                    16'h6FF2: data_out = 8'h83;
                    16'h6FF3: data_out = 8'h84;
                    16'h6FF4: data_out = 8'h85;
                    16'h6FF5: data_out = 8'h86;
                    16'h6FF6: data_out = 8'h87;
                    16'h6FF7: data_out = 8'h88;
                    16'h6FF8: data_out = 8'h89;
                    16'h6FF9: data_out = 8'h8A;
                    16'h6FFA: data_out = 8'h8B;
                    16'h6FFB: data_out = 8'h8C;
                    16'h6FFC: data_out = 8'h8D;
                    16'h6FFD: data_out = 8'h8E;
                    16'h6FFE: data_out = 8'h8F;
                    16'h6FFF: data_out = 8'h90;
                    16'h7000: data_out = 8'h70;
                    16'h7001: data_out = 8'h71;
                    16'h7002: data_out = 8'h72;
                    16'h7003: data_out = 8'h73;
                    16'h7004: data_out = 8'h74;
                    16'h7005: data_out = 8'h75;
                    16'h7006: data_out = 8'h76;
                    16'h7007: data_out = 8'h77;
                    16'h7008: data_out = 8'h78;
                    16'h7009: data_out = 8'h79;
                    16'h700A: data_out = 8'h7A;
                    16'h700B: data_out = 8'h7B;
                    16'h700C: data_out = 8'h7C;
                    16'h700D: data_out = 8'h7D;
                    16'h700E: data_out = 8'h7E;
                    16'h700F: data_out = 8'h7F;
                    16'h7010: data_out = 8'h80;
                    16'h7011: data_out = 8'h81;
                    16'h7012: data_out = 8'h82;
                    16'h7013: data_out = 8'h83;
                    16'h7014: data_out = 8'h84;
                    16'h7015: data_out = 8'h85;
                    16'h7016: data_out = 8'h86;
                    16'h7017: data_out = 8'h87;
                    16'h7018: data_out = 8'h88;
                    16'h7019: data_out = 8'h89;
                    16'h701A: data_out = 8'h8A;
                    16'h701B: data_out = 8'h8B;
                    16'h701C: data_out = 8'h8C;
                    16'h701D: data_out = 8'h8D;
                    16'h701E: data_out = 8'h8E;
                    16'h701F: data_out = 8'h8F;
                    16'h7020: data_out = 8'h90;
                    16'h7021: data_out = 8'h91;
                    16'h7022: data_out = 8'h92;
                    16'h7023: data_out = 8'h93;
                    16'h7024: data_out = 8'h94;
                    16'h7025: data_out = 8'h95;
                    16'h7026: data_out = 8'h96;
                    16'h7027: data_out = 8'h97;
                    16'h7028: data_out = 8'h98;
                    16'h7029: data_out = 8'h99;
                    16'h702A: data_out = 8'h9A;
                    16'h702B: data_out = 8'h9B;
                    16'h702C: data_out = 8'h9C;
                    16'h702D: data_out = 8'h9D;
                    16'h702E: data_out = 8'h9E;
                    16'h702F: data_out = 8'h9F;
                    16'h7030: data_out = 8'hA0;
                    16'h7031: data_out = 8'hA1;
                    16'h7032: data_out = 8'hA2;
                    16'h7033: data_out = 8'hA3;
                    16'h7034: data_out = 8'hA4;
                    16'h7035: data_out = 8'hA5;
                    16'h7036: data_out = 8'hA6;
                    16'h7037: data_out = 8'hA7;
                    16'h7038: data_out = 8'hA8;
                    16'h7039: data_out = 8'hA9;
                    16'h703A: data_out = 8'hAA;
                    16'h703B: data_out = 8'hAB;
                    16'h703C: data_out = 8'hAC;
                    16'h703D: data_out = 8'hAD;
                    16'h703E: data_out = 8'hAE;
                    16'h703F: data_out = 8'hAF;
                    16'h7040: data_out = 8'hB0;
                    16'h7041: data_out = 8'hB1;
                    16'h7042: data_out = 8'hB2;
                    16'h7043: data_out = 8'hB3;
                    16'h7044: data_out = 8'hB4;
                    16'h7045: data_out = 8'hB5;
                    16'h7046: data_out = 8'hB6;
                    16'h7047: data_out = 8'hB7;
                    16'h7048: data_out = 8'hB8;
                    16'h7049: data_out = 8'hB9;
                    16'h704A: data_out = 8'hBA;
                    16'h704B: data_out = 8'hBB;
                    16'h704C: data_out = 8'hBC;
                    16'h704D: data_out = 8'hBD;
                    16'h704E: data_out = 8'hBE;
                    16'h704F: data_out = 8'hBF;
                    16'h7050: data_out = 8'hC0;
                    16'h7051: data_out = 8'hC1;
                    16'h7052: data_out = 8'hC2;
                    16'h7053: data_out = 8'hC3;
                    16'h7054: data_out = 8'hC4;
                    16'h7055: data_out = 8'hC5;
                    16'h7056: data_out = 8'hC6;
                    16'h7057: data_out = 8'hC7;
                    16'h7058: data_out = 8'hC8;
                    16'h7059: data_out = 8'hC9;
                    16'h705A: data_out = 8'hCA;
                    16'h705B: data_out = 8'hCB;
                    16'h705C: data_out = 8'hCC;
                    16'h705D: data_out = 8'hCD;
                    16'h705E: data_out = 8'hCE;
                    16'h705F: data_out = 8'hCF;
                    16'h7060: data_out = 8'hD0;
                    16'h7061: data_out = 8'hD1;
                    16'h7062: data_out = 8'hD2;
                    16'h7063: data_out = 8'hD3;
                    16'h7064: data_out = 8'hD4;
                    16'h7065: data_out = 8'hD5;
                    16'h7066: data_out = 8'hD6;
                    16'h7067: data_out = 8'hD7;
                    16'h7068: data_out = 8'hD8;
                    16'h7069: data_out = 8'hD9;
                    16'h706A: data_out = 8'hDA;
                    16'h706B: data_out = 8'hDB;
                    16'h706C: data_out = 8'hDC;
                    16'h706D: data_out = 8'hDD;
                    16'h706E: data_out = 8'hDE;
                    16'h706F: data_out = 8'hDF;
                    16'h7070: data_out = 8'hE0;
                    16'h7071: data_out = 8'hE1;
                    16'h7072: data_out = 8'hE2;
                    16'h7073: data_out = 8'hE3;
                    16'h7074: data_out = 8'hE4;
                    16'h7075: data_out = 8'hE5;
                    16'h7076: data_out = 8'hE6;
                    16'h7077: data_out = 8'hE7;
                    16'h7078: data_out = 8'hE8;
                    16'h7079: data_out = 8'hE9;
                    16'h707A: data_out = 8'hEA;
                    16'h707B: data_out = 8'hEB;
                    16'h707C: data_out = 8'hEC;
                    16'h707D: data_out = 8'hED;
                    16'h707E: data_out = 8'hEE;
                    16'h707F: data_out = 8'hEF;
                    16'h7080: data_out = 8'h70;
                    16'h7081: data_out = 8'h6F;
                    16'h7082: data_out = 8'h6E;
                    16'h7083: data_out = 8'h6D;
                    16'h7084: data_out = 8'h6C;
                    16'h7085: data_out = 8'h6B;
                    16'h7086: data_out = 8'h6A;
                    16'h7087: data_out = 8'h69;
                    16'h7088: data_out = 8'h68;
                    16'h7089: data_out = 8'h67;
                    16'h708A: data_out = 8'h66;
                    16'h708B: data_out = 8'h65;
                    16'h708C: data_out = 8'h64;
                    16'h708D: data_out = 8'h63;
                    16'h708E: data_out = 8'h62;
                    16'h708F: data_out = 8'h61;
                    16'h7090: data_out = 8'h60;
                    16'h7091: data_out = 8'h5F;
                    16'h7092: data_out = 8'h5E;
                    16'h7093: data_out = 8'h5D;
                    16'h7094: data_out = 8'h5C;
                    16'h7095: data_out = 8'h5B;
                    16'h7096: data_out = 8'h5A;
                    16'h7097: data_out = 8'h59;
                    16'h7098: data_out = 8'h58;
                    16'h7099: data_out = 8'h57;
                    16'h709A: data_out = 8'h56;
                    16'h709B: data_out = 8'h55;
                    16'h709C: data_out = 8'h54;
                    16'h709D: data_out = 8'h53;
                    16'h709E: data_out = 8'h52;
                    16'h709F: data_out = 8'h51;
                    16'h70A0: data_out = 8'h50;
                    16'h70A1: data_out = 8'h4F;
                    16'h70A2: data_out = 8'h4E;
                    16'h70A3: data_out = 8'h4D;
                    16'h70A4: data_out = 8'h4C;
                    16'h70A5: data_out = 8'h4B;
                    16'h70A6: data_out = 8'h4A;
                    16'h70A7: data_out = 8'h49;
                    16'h70A8: data_out = 8'h48;
                    16'h70A9: data_out = 8'h47;
                    16'h70AA: data_out = 8'h46;
                    16'h70AB: data_out = 8'h45;
                    16'h70AC: data_out = 8'h44;
                    16'h70AD: data_out = 8'h43;
                    16'h70AE: data_out = 8'h42;
                    16'h70AF: data_out = 8'h41;
                    16'h70B0: data_out = 8'h40;
                    16'h70B1: data_out = 8'h3F;
                    16'h70B2: data_out = 8'h3E;
                    16'h70B3: data_out = 8'h3D;
                    16'h70B4: data_out = 8'h3C;
                    16'h70B5: data_out = 8'h3B;
                    16'h70B6: data_out = 8'h3A;
                    16'h70B7: data_out = 8'h39;
                    16'h70B8: data_out = 8'h38;
                    16'h70B9: data_out = 8'h37;
                    16'h70BA: data_out = 8'h36;
                    16'h70BB: data_out = 8'h35;
                    16'h70BC: data_out = 8'h34;
                    16'h70BD: data_out = 8'h33;
                    16'h70BE: data_out = 8'h32;
                    16'h70BF: data_out = 8'h31;
                    16'h70C0: data_out = 8'h30;
                    16'h70C1: data_out = 8'h2F;
                    16'h70C2: data_out = 8'h2E;
                    16'h70C3: data_out = 8'h2D;
                    16'h70C4: data_out = 8'h2C;
                    16'h70C5: data_out = 8'h2B;
                    16'h70C6: data_out = 8'h2A;
                    16'h70C7: data_out = 8'h29;
                    16'h70C8: data_out = 8'h28;
                    16'h70C9: data_out = 8'h27;
                    16'h70CA: data_out = 8'h26;
                    16'h70CB: data_out = 8'h25;
                    16'h70CC: data_out = 8'h24;
                    16'h70CD: data_out = 8'h23;
                    16'h70CE: data_out = 8'h22;
                    16'h70CF: data_out = 8'h21;
                    16'h70D0: data_out = 8'h20;
                    16'h70D1: data_out = 8'h1F;
                    16'h70D2: data_out = 8'h1E;
                    16'h70D3: data_out = 8'h1D;
                    16'h70D4: data_out = 8'h1C;
                    16'h70D5: data_out = 8'h1B;
                    16'h70D6: data_out = 8'h1A;
                    16'h70D7: data_out = 8'h19;
                    16'h70D8: data_out = 8'h18;
                    16'h70D9: data_out = 8'h17;
                    16'h70DA: data_out = 8'h16;
                    16'h70DB: data_out = 8'h15;
                    16'h70DC: data_out = 8'h14;
                    16'h70DD: data_out = 8'h13;
                    16'h70DE: data_out = 8'h12;
                    16'h70DF: data_out = 8'h11;
                    16'h70E0: data_out = 8'h10;
                    16'h70E1: data_out = 8'hF;
                    16'h70E2: data_out = 8'hE;
                    16'h70E3: data_out = 8'hD;
                    16'h70E4: data_out = 8'hC;
                    16'h70E5: data_out = 8'hB;
                    16'h70E6: data_out = 8'hA;
                    16'h70E7: data_out = 8'h9;
                    16'h70E8: data_out = 8'h8;
                    16'h70E9: data_out = 8'h7;
                    16'h70EA: data_out = 8'h6;
                    16'h70EB: data_out = 8'h5;
                    16'h70EC: data_out = 8'h4;
                    16'h70ED: data_out = 8'h3;
                    16'h70EE: data_out = 8'h2;
                    16'h70EF: data_out = 8'h1;
                    16'h70F0: data_out = 8'h0;
                    16'h70F1: data_out = 8'h81;
                    16'h70F2: data_out = 8'h82;
                    16'h70F3: data_out = 8'h83;
                    16'h70F4: data_out = 8'h84;
                    16'h70F5: data_out = 8'h85;
                    16'h70F6: data_out = 8'h86;
                    16'h70F7: data_out = 8'h87;
                    16'h70F8: data_out = 8'h88;
                    16'h70F9: data_out = 8'h89;
                    16'h70FA: data_out = 8'h8A;
                    16'h70FB: data_out = 8'h8B;
                    16'h70FC: data_out = 8'h8C;
                    16'h70FD: data_out = 8'h8D;
                    16'h70FE: data_out = 8'h8E;
                    16'h70FF: data_out = 8'h8F;
                    16'h7100: data_out = 8'h71;
                    16'h7101: data_out = 8'h72;
                    16'h7102: data_out = 8'h73;
                    16'h7103: data_out = 8'h74;
                    16'h7104: data_out = 8'h75;
                    16'h7105: data_out = 8'h76;
                    16'h7106: data_out = 8'h77;
                    16'h7107: data_out = 8'h78;
                    16'h7108: data_out = 8'h79;
                    16'h7109: data_out = 8'h7A;
                    16'h710A: data_out = 8'h7B;
                    16'h710B: data_out = 8'h7C;
                    16'h710C: data_out = 8'h7D;
                    16'h710D: data_out = 8'h7E;
                    16'h710E: data_out = 8'h7F;
                    16'h710F: data_out = 8'h80;
                    16'h7110: data_out = 8'h81;
                    16'h7111: data_out = 8'h82;
                    16'h7112: data_out = 8'h83;
                    16'h7113: data_out = 8'h84;
                    16'h7114: data_out = 8'h85;
                    16'h7115: data_out = 8'h86;
                    16'h7116: data_out = 8'h87;
                    16'h7117: data_out = 8'h88;
                    16'h7118: data_out = 8'h89;
                    16'h7119: data_out = 8'h8A;
                    16'h711A: data_out = 8'h8B;
                    16'h711B: data_out = 8'h8C;
                    16'h711C: data_out = 8'h8D;
                    16'h711D: data_out = 8'h8E;
                    16'h711E: data_out = 8'h8F;
                    16'h711F: data_out = 8'h90;
                    16'h7120: data_out = 8'h91;
                    16'h7121: data_out = 8'h92;
                    16'h7122: data_out = 8'h93;
                    16'h7123: data_out = 8'h94;
                    16'h7124: data_out = 8'h95;
                    16'h7125: data_out = 8'h96;
                    16'h7126: data_out = 8'h97;
                    16'h7127: data_out = 8'h98;
                    16'h7128: data_out = 8'h99;
                    16'h7129: data_out = 8'h9A;
                    16'h712A: data_out = 8'h9B;
                    16'h712B: data_out = 8'h9C;
                    16'h712C: data_out = 8'h9D;
                    16'h712D: data_out = 8'h9E;
                    16'h712E: data_out = 8'h9F;
                    16'h712F: data_out = 8'hA0;
                    16'h7130: data_out = 8'hA1;
                    16'h7131: data_out = 8'hA2;
                    16'h7132: data_out = 8'hA3;
                    16'h7133: data_out = 8'hA4;
                    16'h7134: data_out = 8'hA5;
                    16'h7135: data_out = 8'hA6;
                    16'h7136: data_out = 8'hA7;
                    16'h7137: data_out = 8'hA8;
                    16'h7138: data_out = 8'hA9;
                    16'h7139: data_out = 8'hAA;
                    16'h713A: data_out = 8'hAB;
                    16'h713B: data_out = 8'hAC;
                    16'h713C: data_out = 8'hAD;
                    16'h713D: data_out = 8'hAE;
                    16'h713E: data_out = 8'hAF;
                    16'h713F: data_out = 8'hB0;
                    16'h7140: data_out = 8'hB1;
                    16'h7141: data_out = 8'hB2;
                    16'h7142: data_out = 8'hB3;
                    16'h7143: data_out = 8'hB4;
                    16'h7144: data_out = 8'hB5;
                    16'h7145: data_out = 8'hB6;
                    16'h7146: data_out = 8'hB7;
                    16'h7147: data_out = 8'hB8;
                    16'h7148: data_out = 8'hB9;
                    16'h7149: data_out = 8'hBA;
                    16'h714A: data_out = 8'hBB;
                    16'h714B: data_out = 8'hBC;
                    16'h714C: data_out = 8'hBD;
                    16'h714D: data_out = 8'hBE;
                    16'h714E: data_out = 8'hBF;
                    16'h714F: data_out = 8'hC0;
                    16'h7150: data_out = 8'hC1;
                    16'h7151: data_out = 8'hC2;
                    16'h7152: data_out = 8'hC3;
                    16'h7153: data_out = 8'hC4;
                    16'h7154: data_out = 8'hC5;
                    16'h7155: data_out = 8'hC6;
                    16'h7156: data_out = 8'hC7;
                    16'h7157: data_out = 8'hC8;
                    16'h7158: data_out = 8'hC9;
                    16'h7159: data_out = 8'hCA;
                    16'h715A: data_out = 8'hCB;
                    16'h715B: data_out = 8'hCC;
                    16'h715C: data_out = 8'hCD;
                    16'h715D: data_out = 8'hCE;
                    16'h715E: data_out = 8'hCF;
                    16'h715F: data_out = 8'hD0;
                    16'h7160: data_out = 8'hD1;
                    16'h7161: data_out = 8'hD2;
                    16'h7162: data_out = 8'hD3;
                    16'h7163: data_out = 8'hD4;
                    16'h7164: data_out = 8'hD5;
                    16'h7165: data_out = 8'hD6;
                    16'h7166: data_out = 8'hD7;
                    16'h7167: data_out = 8'hD8;
                    16'h7168: data_out = 8'hD9;
                    16'h7169: data_out = 8'hDA;
                    16'h716A: data_out = 8'hDB;
                    16'h716B: data_out = 8'hDC;
                    16'h716C: data_out = 8'hDD;
                    16'h716D: data_out = 8'hDE;
                    16'h716E: data_out = 8'hDF;
                    16'h716F: data_out = 8'hE0;
                    16'h7170: data_out = 8'hE1;
                    16'h7171: data_out = 8'hE2;
                    16'h7172: data_out = 8'hE3;
                    16'h7173: data_out = 8'hE4;
                    16'h7174: data_out = 8'hE5;
                    16'h7175: data_out = 8'hE6;
                    16'h7176: data_out = 8'hE7;
                    16'h7177: data_out = 8'hE8;
                    16'h7178: data_out = 8'hE9;
                    16'h7179: data_out = 8'hEA;
                    16'h717A: data_out = 8'hEB;
                    16'h717B: data_out = 8'hEC;
                    16'h717C: data_out = 8'hED;
                    16'h717D: data_out = 8'hEE;
                    16'h717E: data_out = 8'hEF;
                    16'h717F: data_out = 8'hF0;
                    16'h7180: data_out = 8'h71;
                    16'h7181: data_out = 8'h70;
                    16'h7182: data_out = 8'h6F;
                    16'h7183: data_out = 8'h6E;
                    16'h7184: data_out = 8'h6D;
                    16'h7185: data_out = 8'h6C;
                    16'h7186: data_out = 8'h6B;
                    16'h7187: data_out = 8'h6A;
                    16'h7188: data_out = 8'h69;
                    16'h7189: data_out = 8'h68;
                    16'h718A: data_out = 8'h67;
                    16'h718B: data_out = 8'h66;
                    16'h718C: data_out = 8'h65;
                    16'h718D: data_out = 8'h64;
                    16'h718E: data_out = 8'h63;
                    16'h718F: data_out = 8'h62;
                    16'h7190: data_out = 8'h61;
                    16'h7191: data_out = 8'h60;
                    16'h7192: data_out = 8'h5F;
                    16'h7193: data_out = 8'h5E;
                    16'h7194: data_out = 8'h5D;
                    16'h7195: data_out = 8'h5C;
                    16'h7196: data_out = 8'h5B;
                    16'h7197: data_out = 8'h5A;
                    16'h7198: data_out = 8'h59;
                    16'h7199: data_out = 8'h58;
                    16'h719A: data_out = 8'h57;
                    16'h719B: data_out = 8'h56;
                    16'h719C: data_out = 8'h55;
                    16'h719D: data_out = 8'h54;
                    16'h719E: data_out = 8'h53;
                    16'h719F: data_out = 8'h52;
                    16'h71A0: data_out = 8'h51;
                    16'h71A1: data_out = 8'h50;
                    16'h71A2: data_out = 8'h4F;
                    16'h71A3: data_out = 8'h4E;
                    16'h71A4: data_out = 8'h4D;
                    16'h71A5: data_out = 8'h4C;
                    16'h71A6: data_out = 8'h4B;
                    16'h71A7: data_out = 8'h4A;
                    16'h71A8: data_out = 8'h49;
                    16'h71A9: data_out = 8'h48;
                    16'h71AA: data_out = 8'h47;
                    16'h71AB: data_out = 8'h46;
                    16'h71AC: data_out = 8'h45;
                    16'h71AD: data_out = 8'h44;
                    16'h71AE: data_out = 8'h43;
                    16'h71AF: data_out = 8'h42;
                    16'h71B0: data_out = 8'h41;
                    16'h71B1: data_out = 8'h40;
                    16'h71B2: data_out = 8'h3F;
                    16'h71B3: data_out = 8'h3E;
                    16'h71B4: data_out = 8'h3D;
                    16'h71B5: data_out = 8'h3C;
                    16'h71B6: data_out = 8'h3B;
                    16'h71B7: data_out = 8'h3A;
                    16'h71B8: data_out = 8'h39;
                    16'h71B9: data_out = 8'h38;
                    16'h71BA: data_out = 8'h37;
                    16'h71BB: data_out = 8'h36;
                    16'h71BC: data_out = 8'h35;
                    16'h71BD: data_out = 8'h34;
                    16'h71BE: data_out = 8'h33;
                    16'h71BF: data_out = 8'h32;
                    16'h71C0: data_out = 8'h31;
                    16'h71C1: data_out = 8'h30;
                    16'h71C2: data_out = 8'h2F;
                    16'h71C3: data_out = 8'h2E;
                    16'h71C4: data_out = 8'h2D;
                    16'h71C5: data_out = 8'h2C;
                    16'h71C6: data_out = 8'h2B;
                    16'h71C7: data_out = 8'h2A;
                    16'h71C8: data_out = 8'h29;
                    16'h71C9: data_out = 8'h28;
                    16'h71CA: data_out = 8'h27;
                    16'h71CB: data_out = 8'h26;
                    16'h71CC: data_out = 8'h25;
                    16'h71CD: data_out = 8'h24;
                    16'h71CE: data_out = 8'h23;
                    16'h71CF: data_out = 8'h22;
                    16'h71D0: data_out = 8'h21;
                    16'h71D1: data_out = 8'h20;
                    16'h71D2: data_out = 8'h1F;
                    16'h71D3: data_out = 8'h1E;
                    16'h71D4: data_out = 8'h1D;
                    16'h71D5: data_out = 8'h1C;
                    16'h71D6: data_out = 8'h1B;
                    16'h71D7: data_out = 8'h1A;
                    16'h71D8: data_out = 8'h19;
                    16'h71D9: data_out = 8'h18;
                    16'h71DA: data_out = 8'h17;
                    16'h71DB: data_out = 8'h16;
                    16'h71DC: data_out = 8'h15;
                    16'h71DD: data_out = 8'h14;
                    16'h71DE: data_out = 8'h13;
                    16'h71DF: data_out = 8'h12;
                    16'h71E0: data_out = 8'h11;
                    16'h71E1: data_out = 8'h10;
                    16'h71E2: data_out = 8'hF;
                    16'h71E3: data_out = 8'hE;
                    16'h71E4: data_out = 8'hD;
                    16'h71E5: data_out = 8'hC;
                    16'h71E6: data_out = 8'hB;
                    16'h71E7: data_out = 8'hA;
                    16'h71E8: data_out = 8'h9;
                    16'h71E9: data_out = 8'h8;
                    16'h71EA: data_out = 8'h7;
                    16'h71EB: data_out = 8'h6;
                    16'h71EC: data_out = 8'h5;
                    16'h71ED: data_out = 8'h4;
                    16'h71EE: data_out = 8'h3;
                    16'h71EF: data_out = 8'h2;
                    16'h71F0: data_out = 8'h1;
                    16'h71F1: data_out = 8'h0;
                    16'h71F2: data_out = 8'h81;
                    16'h71F3: data_out = 8'h82;
                    16'h71F4: data_out = 8'h83;
                    16'h71F5: data_out = 8'h84;
                    16'h71F6: data_out = 8'h85;
                    16'h71F7: data_out = 8'h86;
                    16'h71F8: data_out = 8'h87;
                    16'h71F9: data_out = 8'h88;
                    16'h71FA: data_out = 8'h89;
                    16'h71FB: data_out = 8'h8A;
                    16'h71FC: data_out = 8'h8B;
                    16'h71FD: data_out = 8'h8C;
                    16'h71FE: data_out = 8'h8D;
                    16'h71FF: data_out = 8'h8E;
                    16'h7200: data_out = 8'h72;
                    16'h7201: data_out = 8'h73;
                    16'h7202: data_out = 8'h74;
                    16'h7203: data_out = 8'h75;
                    16'h7204: data_out = 8'h76;
                    16'h7205: data_out = 8'h77;
                    16'h7206: data_out = 8'h78;
                    16'h7207: data_out = 8'h79;
                    16'h7208: data_out = 8'h7A;
                    16'h7209: data_out = 8'h7B;
                    16'h720A: data_out = 8'h7C;
                    16'h720B: data_out = 8'h7D;
                    16'h720C: data_out = 8'h7E;
                    16'h720D: data_out = 8'h7F;
                    16'h720E: data_out = 8'h80;
                    16'h720F: data_out = 8'h81;
                    16'h7210: data_out = 8'h82;
                    16'h7211: data_out = 8'h83;
                    16'h7212: data_out = 8'h84;
                    16'h7213: data_out = 8'h85;
                    16'h7214: data_out = 8'h86;
                    16'h7215: data_out = 8'h87;
                    16'h7216: data_out = 8'h88;
                    16'h7217: data_out = 8'h89;
                    16'h7218: data_out = 8'h8A;
                    16'h7219: data_out = 8'h8B;
                    16'h721A: data_out = 8'h8C;
                    16'h721B: data_out = 8'h8D;
                    16'h721C: data_out = 8'h8E;
                    16'h721D: data_out = 8'h8F;
                    16'h721E: data_out = 8'h90;
                    16'h721F: data_out = 8'h91;
                    16'h7220: data_out = 8'h92;
                    16'h7221: data_out = 8'h93;
                    16'h7222: data_out = 8'h94;
                    16'h7223: data_out = 8'h95;
                    16'h7224: data_out = 8'h96;
                    16'h7225: data_out = 8'h97;
                    16'h7226: data_out = 8'h98;
                    16'h7227: data_out = 8'h99;
                    16'h7228: data_out = 8'h9A;
                    16'h7229: data_out = 8'h9B;
                    16'h722A: data_out = 8'h9C;
                    16'h722B: data_out = 8'h9D;
                    16'h722C: data_out = 8'h9E;
                    16'h722D: data_out = 8'h9F;
                    16'h722E: data_out = 8'hA0;
                    16'h722F: data_out = 8'hA1;
                    16'h7230: data_out = 8'hA2;
                    16'h7231: data_out = 8'hA3;
                    16'h7232: data_out = 8'hA4;
                    16'h7233: data_out = 8'hA5;
                    16'h7234: data_out = 8'hA6;
                    16'h7235: data_out = 8'hA7;
                    16'h7236: data_out = 8'hA8;
                    16'h7237: data_out = 8'hA9;
                    16'h7238: data_out = 8'hAA;
                    16'h7239: data_out = 8'hAB;
                    16'h723A: data_out = 8'hAC;
                    16'h723B: data_out = 8'hAD;
                    16'h723C: data_out = 8'hAE;
                    16'h723D: data_out = 8'hAF;
                    16'h723E: data_out = 8'hB0;
                    16'h723F: data_out = 8'hB1;
                    16'h7240: data_out = 8'hB2;
                    16'h7241: data_out = 8'hB3;
                    16'h7242: data_out = 8'hB4;
                    16'h7243: data_out = 8'hB5;
                    16'h7244: data_out = 8'hB6;
                    16'h7245: data_out = 8'hB7;
                    16'h7246: data_out = 8'hB8;
                    16'h7247: data_out = 8'hB9;
                    16'h7248: data_out = 8'hBA;
                    16'h7249: data_out = 8'hBB;
                    16'h724A: data_out = 8'hBC;
                    16'h724B: data_out = 8'hBD;
                    16'h724C: data_out = 8'hBE;
                    16'h724D: data_out = 8'hBF;
                    16'h724E: data_out = 8'hC0;
                    16'h724F: data_out = 8'hC1;
                    16'h7250: data_out = 8'hC2;
                    16'h7251: data_out = 8'hC3;
                    16'h7252: data_out = 8'hC4;
                    16'h7253: data_out = 8'hC5;
                    16'h7254: data_out = 8'hC6;
                    16'h7255: data_out = 8'hC7;
                    16'h7256: data_out = 8'hC8;
                    16'h7257: data_out = 8'hC9;
                    16'h7258: data_out = 8'hCA;
                    16'h7259: data_out = 8'hCB;
                    16'h725A: data_out = 8'hCC;
                    16'h725B: data_out = 8'hCD;
                    16'h725C: data_out = 8'hCE;
                    16'h725D: data_out = 8'hCF;
                    16'h725E: data_out = 8'hD0;
                    16'h725F: data_out = 8'hD1;
                    16'h7260: data_out = 8'hD2;
                    16'h7261: data_out = 8'hD3;
                    16'h7262: data_out = 8'hD4;
                    16'h7263: data_out = 8'hD5;
                    16'h7264: data_out = 8'hD6;
                    16'h7265: data_out = 8'hD7;
                    16'h7266: data_out = 8'hD8;
                    16'h7267: data_out = 8'hD9;
                    16'h7268: data_out = 8'hDA;
                    16'h7269: data_out = 8'hDB;
                    16'h726A: data_out = 8'hDC;
                    16'h726B: data_out = 8'hDD;
                    16'h726C: data_out = 8'hDE;
                    16'h726D: data_out = 8'hDF;
                    16'h726E: data_out = 8'hE0;
                    16'h726F: data_out = 8'hE1;
                    16'h7270: data_out = 8'hE2;
                    16'h7271: data_out = 8'hE3;
                    16'h7272: data_out = 8'hE4;
                    16'h7273: data_out = 8'hE5;
                    16'h7274: data_out = 8'hE6;
                    16'h7275: data_out = 8'hE7;
                    16'h7276: data_out = 8'hE8;
                    16'h7277: data_out = 8'hE9;
                    16'h7278: data_out = 8'hEA;
                    16'h7279: data_out = 8'hEB;
                    16'h727A: data_out = 8'hEC;
                    16'h727B: data_out = 8'hED;
                    16'h727C: data_out = 8'hEE;
                    16'h727D: data_out = 8'hEF;
                    16'h727E: data_out = 8'hF0;
                    16'h727F: data_out = 8'hF1;
                    16'h7280: data_out = 8'h72;
                    16'h7281: data_out = 8'h71;
                    16'h7282: data_out = 8'h70;
                    16'h7283: data_out = 8'h6F;
                    16'h7284: data_out = 8'h6E;
                    16'h7285: data_out = 8'h6D;
                    16'h7286: data_out = 8'h6C;
                    16'h7287: data_out = 8'h6B;
                    16'h7288: data_out = 8'h6A;
                    16'h7289: data_out = 8'h69;
                    16'h728A: data_out = 8'h68;
                    16'h728B: data_out = 8'h67;
                    16'h728C: data_out = 8'h66;
                    16'h728D: data_out = 8'h65;
                    16'h728E: data_out = 8'h64;
                    16'h728F: data_out = 8'h63;
                    16'h7290: data_out = 8'h62;
                    16'h7291: data_out = 8'h61;
                    16'h7292: data_out = 8'h60;
                    16'h7293: data_out = 8'h5F;
                    16'h7294: data_out = 8'h5E;
                    16'h7295: data_out = 8'h5D;
                    16'h7296: data_out = 8'h5C;
                    16'h7297: data_out = 8'h5B;
                    16'h7298: data_out = 8'h5A;
                    16'h7299: data_out = 8'h59;
                    16'h729A: data_out = 8'h58;
                    16'h729B: data_out = 8'h57;
                    16'h729C: data_out = 8'h56;
                    16'h729D: data_out = 8'h55;
                    16'h729E: data_out = 8'h54;
                    16'h729F: data_out = 8'h53;
                    16'h72A0: data_out = 8'h52;
                    16'h72A1: data_out = 8'h51;
                    16'h72A2: data_out = 8'h50;
                    16'h72A3: data_out = 8'h4F;
                    16'h72A4: data_out = 8'h4E;
                    16'h72A5: data_out = 8'h4D;
                    16'h72A6: data_out = 8'h4C;
                    16'h72A7: data_out = 8'h4B;
                    16'h72A8: data_out = 8'h4A;
                    16'h72A9: data_out = 8'h49;
                    16'h72AA: data_out = 8'h48;
                    16'h72AB: data_out = 8'h47;
                    16'h72AC: data_out = 8'h46;
                    16'h72AD: data_out = 8'h45;
                    16'h72AE: data_out = 8'h44;
                    16'h72AF: data_out = 8'h43;
                    16'h72B0: data_out = 8'h42;
                    16'h72B1: data_out = 8'h41;
                    16'h72B2: data_out = 8'h40;
                    16'h72B3: data_out = 8'h3F;
                    16'h72B4: data_out = 8'h3E;
                    16'h72B5: data_out = 8'h3D;
                    16'h72B6: data_out = 8'h3C;
                    16'h72B7: data_out = 8'h3B;
                    16'h72B8: data_out = 8'h3A;
                    16'h72B9: data_out = 8'h39;
                    16'h72BA: data_out = 8'h38;
                    16'h72BB: data_out = 8'h37;
                    16'h72BC: data_out = 8'h36;
                    16'h72BD: data_out = 8'h35;
                    16'h72BE: data_out = 8'h34;
                    16'h72BF: data_out = 8'h33;
                    16'h72C0: data_out = 8'h32;
                    16'h72C1: data_out = 8'h31;
                    16'h72C2: data_out = 8'h30;
                    16'h72C3: data_out = 8'h2F;
                    16'h72C4: data_out = 8'h2E;
                    16'h72C5: data_out = 8'h2D;
                    16'h72C6: data_out = 8'h2C;
                    16'h72C7: data_out = 8'h2B;
                    16'h72C8: data_out = 8'h2A;
                    16'h72C9: data_out = 8'h29;
                    16'h72CA: data_out = 8'h28;
                    16'h72CB: data_out = 8'h27;
                    16'h72CC: data_out = 8'h26;
                    16'h72CD: data_out = 8'h25;
                    16'h72CE: data_out = 8'h24;
                    16'h72CF: data_out = 8'h23;
                    16'h72D0: data_out = 8'h22;
                    16'h72D1: data_out = 8'h21;
                    16'h72D2: data_out = 8'h20;
                    16'h72D3: data_out = 8'h1F;
                    16'h72D4: data_out = 8'h1E;
                    16'h72D5: data_out = 8'h1D;
                    16'h72D6: data_out = 8'h1C;
                    16'h72D7: data_out = 8'h1B;
                    16'h72D8: data_out = 8'h1A;
                    16'h72D9: data_out = 8'h19;
                    16'h72DA: data_out = 8'h18;
                    16'h72DB: data_out = 8'h17;
                    16'h72DC: data_out = 8'h16;
                    16'h72DD: data_out = 8'h15;
                    16'h72DE: data_out = 8'h14;
                    16'h72DF: data_out = 8'h13;
                    16'h72E0: data_out = 8'h12;
                    16'h72E1: data_out = 8'h11;
                    16'h72E2: data_out = 8'h10;
                    16'h72E3: data_out = 8'hF;
                    16'h72E4: data_out = 8'hE;
                    16'h72E5: data_out = 8'hD;
                    16'h72E6: data_out = 8'hC;
                    16'h72E7: data_out = 8'hB;
                    16'h72E8: data_out = 8'hA;
                    16'h72E9: data_out = 8'h9;
                    16'h72EA: data_out = 8'h8;
                    16'h72EB: data_out = 8'h7;
                    16'h72EC: data_out = 8'h6;
                    16'h72ED: data_out = 8'h5;
                    16'h72EE: data_out = 8'h4;
                    16'h72EF: data_out = 8'h3;
                    16'h72F0: data_out = 8'h2;
                    16'h72F1: data_out = 8'h1;
                    16'h72F2: data_out = 8'h0;
                    16'h72F3: data_out = 8'h81;
                    16'h72F4: data_out = 8'h82;
                    16'h72F5: data_out = 8'h83;
                    16'h72F6: data_out = 8'h84;
                    16'h72F7: data_out = 8'h85;
                    16'h72F8: data_out = 8'h86;
                    16'h72F9: data_out = 8'h87;
                    16'h72FA: data_out = 8'h88;
                    16'h72FB: data_out = 8'h89;
                    16'h72FC: data_out = 8'h8A;
                    16'h72FD: data_out = 8'h8B;
                    16'h72FE: data_out = 8'h8C;
                    16'h72FF: data_out = 8'h8D;
                    16'h7300: data_out = 8'h73;
                    16'h7301: data_out = 8'h74;
                    16'h7302: data_out = 8'h75;
                    16'h7303: data_out = 8'h76;
                    16'h7304: data_out = 8'h77;
                    16'h7305: data_out = 8'h78;
                    16'h7306: data_out = 8'h79;
                    16'h7307: data_out = 8'h7A;
                    16'h7308: data_out = 8'h7B;
                    16'h7309: data_out = 8'h7C;
                    16'h730A: data_out = 8'h7D;
                    16'h730B: data_out = 8'h7E;
                    16'h730C: data_out = 8'h7F;
                    16'h730D: data_out = 8'h80;
                    16'h730E: data_out = 8'h81;
                    16'h730F: data_out = 8'h82;
                    16'h7310: data_out = 8'h83;
                    16'h7311: data_out = 8'h84;
                    16'h7312: data_out = 8'h85;
                    16'h7313: data_out = 8'h86;
                    16'h7314: data_out = 8'h87;
                    16'h7315: data_out = 8'h88;
                    16'h7316: data_out = 8'h89;
                    16'h7317: data_out = 8'h8A;
                    16'h7318: data_out = 8'h8B;
                    16'h7319: data_out = 8'h8C;
                    16'h731A: data_out = 8'h8D;
                    16'h731B: data_out = 8'h8E;
                    16'h731C: data_out = 8'h8F;
                    16'h731D: data_out = 8'h90;
                    16'h731E: data_out = 8'h91;
                    16'h731F: data_out = 8'h92;
                    16'h7320: data_out = 8'h93;
                    16'h7321: data_out = 8'h94;
                    16'h7322: data_out = 8'h95;
                    16'h7323: data_out = 8'h96;
                    16'h7324: data_out = 8'h97;
                    16'h7325: data_out = 8'h98;
                    16'h7326: data_out = 8'h99;
                    16'h7327: data_out = 8'h9A;
                    16'h7328: data_out = 8'h9B;
                    16'h7329: data_out = 8'h9C;
                    16'h732A: data_out = 8'h9D;
                    16'h732B: data_out = 8'h9E;
                    16'h732C: data_out = 8'h9F;
                    16'h732D: data_out = 8'hA0;
                    16'h732E: data_out = 8'hA1;
                    16'h732F: data_out = 8'hA2;
                    16'h7330: data_out = 8'hA3;
                    16'h7331: data_out = 8'hA4;
                    16'h7332: data_out = 8'hA5;
                    16'h7333: data_out = 8'hA6;
                    16'h7334: data_out = 8'hA7;
                    16'h7335: data_out = 8'hA8;
                    16'h7336: data_out = 8'hA9;
                    16'h7337: data_out = 8'hAA;
                    16'h7338: data_out = 8'hAB;
                    16'h7339: data_out = 8'hAC;
                    16'h733A: data_out = 8'hAD;
                    16'h733B: data_out = 8'hAE;
                    16'h733C: data_out = 8'hAF;
                    16'h733D: data_out = 8'hB0;
                    16'h733E: data_out = 8'hB1;
                    16'h733F: data_out = 8'hB2;
                    16'h7340: data_out = 8'hB3;
                    16'h7341: data_out = 8'hB4;
                    16'h7342: data_out = 8'hB5;
                    16'h7343: data_out = 8'hB6;
                    16'h7344: data_out = 8'hB7;
                    16'h7345: data_out = 8'hB8;
                    16'h7346: data_out = 8'hB9;
                    16'h7347: data_out = 8'hBA;
                    16'h7348: data_out = 8'hBB;
                    16'h7349: data_out = 8'hBC;
                    16'h734A: data_out = 8'hBD;
                    16'h734B: data_out = 8'hBE;
                    16'h734C: data_out = 8'hBF;
                    16'h734D: data_out = 8'hC0;
                    16'h734E: data_out = 8'hC1;
                    16'h734F: data_out = 8'hC2;
                    16'h7350: data_out = 8'hC3;
                    16'h7351: data_out = 8'hC4;
                    16'h7352: data_out = 8'hC5;
                    16'h7353: data_out = 8'hC6;
                    16'h7354: data_out = 8'hC7;
                    16'h7355: data_out = 8'hC8;
                    16'h7356: data_out = 8'hC9;
                    16'h7357: data_out = 8'hCA;
                    16'h7358: data_out = 8'hCB;
                    16'h7359: data_out = 8'hCC;
                    16'h735A: data_out = 8'hCD;
                    16'h735B: data_out = 8'hCE;
                    16'h735C: data_out = 8'hCF;
                    16'h735D: data_out = 8'hD0;
                    16'h735E: data_out = 8'hD1;
                    16'h735F: data_out = 8'hD2;
                    16'h7360: data_out = 8'hD3;
                    16'h7361: data_out = 8'hD4;
                    16'h7362: data_out = 8'hD5;
                    16'h7363: data_out = 8'hD6;
                    16'h7364: data_out = 8'hD7;
                    16'h7365: data_out = 8'hD8;
                    16'h7366: data_out = 8'hD9;
                    16'h7367: data_out = 8'hDA;
                    16'h7368: data_out = 8'hDB;
                    16'h7369: data_out = 8'hDC;
                    16'h736A: data_out = 8'hDD;
                    16'h736B: data_out = 8'hDE;
                    16'h736C: data_out = 8'hDF;
                    16'h736D: data_out = 8'hE0;
                    16'h736E: data_out = 8'hE1;
                    16'h736F: data_out = 8'hE2;
                    16'h7370: data_out = 8'hE3;
                    16'h7371: data_out = 8'hE4;
                    16'h7372: data_out = 8'hE5;
                    16'h7373: data_out = 8'hE6;
                    16'h7374: data_out = 8'hE7;
                    16'h7375: data_out = 8'hE8;
                    16'h7376: data_out = 8'hE9;
                    16'h7377: data_out = 8'hEA;
                    16'h7378: data_out = 8'hEB;
                    16'h7379: data_out = 8'hEC;
                    16'h737A: data_out = 8'hED;
                    16'h737B: data_out = 8'hEE;
                    16'h737C: data_out = 8'hEF;
                    16'h737D: data_out = 8'hF0;
                    16'h737E: data_out = 8'hF1;
                    16'h737F: data_out = 8'hF2;
                    16'h7380: data_out = 8'h73;
                    16'h7381: data_out = 8'h72;
                    16'h7382: data_out = 8'h71;
                    16'h7383: data_out = 8'h70;
                    16'h7384: data_out = 8'h6F;
                    16'h7385: data_out = 8'h6E;
                    16'h7386: data_out = 8'h6D;
                    16'h7387: data_out = 8'h6C;
                    16'h7388: data_out = 8'h6B;
                    16'h7389: data_out = 8'h6A;
                    16'h738A: data_out = 8'h69;
                    16'h738B: data_out = 8'h68;
                    16'h738C: data_out = 8'h67;
                    16'h738D: data_out = 8'h66;
                    16'h738E: data_out = 8'h65;
                    16'h738F: data_out = 8'h64;
                    16'h7390: data_out = 8'h63;
                    16'h7391: data_out = 8'h62;
                    16'h7392: data_out = 8'h61;
                    16'h7393: data_out = 8'h60;
                    16'h7394: data_out = 8'h5F;
                    16'h7395: data_out = 8'h5E;
                    16'h7396: data_out = 8'h5D;
                    16'h7397: data_out = 8'h5C;
                    16'h7398: data_out = 8'h5B;
                    16'h7399: data_out = 8'h5A;
                    16'h739A: data_out = 8'h59;
                    16'h739B: data_out = 8'h58;
                    16'h739C: data_out = 8'h57;
                    16'h739D: data_out = 8'h56;
                    16'h739E: data_out = 8'h55;
                    16'h739F: data_out = 8'h54;
                    16'h73A0: data_out = 8'h53;
                    16'h73A1: data_out = 8'h52;
                    16'h73A2: data_out = 8'h51;
                    16'h73A3: data_out = 8'h50;
                    16'h73A4: data_out = 8'h4F;
                    16'h73A5: data_out = 8'h4E;
                    16'h73A6: data_out = 8'h4D;
                    16'h73A7: data_out = 8'h4C;
                    16'h73A8: data_out = 8'h4B;
                    16'h73A9: data_out = 8'h4A;
                    16'h73AA: data_out = 8'h49;
                    16'h73AB: data_out = 8'h48;
                    16'h73AC: data_out = 8'h47;
                    16'h73AD: data_out = 8'h46;
                    16'h73AE: data_out = 8'h45;
                    16'h73AF: data_out = 8'h44;
                    16'h73B0: data_out = 8'h43;
                    16'h73B1: data_out = 8'h42;
                    16'h73B2: data_out = 8'h41;
                    16'h73B3: data_out = 8'h40;
                    16'h73B4: data_out = 8'h3F;
                    16'h73B5: data_out = 8'h3E;
                    16'h73B6: data_out = 8'h3D;
                    16'h73B7: data_out = 8'h3C;
                    16'h73B8: data_out = 8'h3B;
                    16'h73B9: data_out = 8'h3A;
                    16'h73BA: data_out = 8'h39;
                    16'h73BB: data_out = 8'h38;
                    16'h73BC: data_out = 8'h37;
                    16'h73BD: data_out = 8'h36;
                    16'h73BE: data_out = 8'h35;
                    16'h73BF: data_out = 8'h34;
                    16'h73C0: data_out = 8'h33;
                    16'h73C1: data_out = 8'h32;
                    16'h73C2: data_out = 8'h31;
                    16'h73C3: data_out = 8'h30;
                    16'h73C4: data_out = 8'h2F;
                    16'h73C5: data_out = 8'h2E;
                    16'h73C6: data_out = 8'h2D;
                    16'h73C7: data_out = 8'h2C;
                    16'h73C8: data_out = 8'h2B;
                    16'h73C9: data_out = 8'h2A;
                    16'h73CA: data_out = 8'h29;
                    16'h73CB: data_out = 8'h28;
                    16'h73CC: data_out = 8'h27;
                    16'h73CD: data_out = 8'h26;
                    16'h73CE: data_out = 8'h25;
                    16'h73CF: data_out = 8'h24;
                    16'h73D0: data_out = 8'h23;
                    16'h73D1: data_out = 8'h22;
                    16'h73D2: data_out = 8'h21;
                    16'h73D3: data_out = 8'h20;
                    16'h73D4: data_out = 8'h1F;
                    16'h73D5: data_out = 8'h1E;
                    16'h73D6: data_out = 8'h1D;
                    16'h73D7: data_out = 8'h1C;
                    16'h73D8: data_out = 8'h1B;
                    16'h73D9: data_out = 8'h1A;
                    16'h73DA: data_out = 8'h19;
                    16'h73DB: data_out = 8'h18;
                    16'h73DC: data_out = 8'h17;
                    16'h73DD: data_out = 8'h16;
                    16'h73DE: data_out = 8'h15;
                    16'h73DF: data_out = 8'h14;
                    16'h73E0: data_out = 8'h13;
                    16'h73E1: data_out = 8'h12;
                    16'h73E2: data_out = 8'h11;
                    16'h73E3: data_out = 8'h10;
                    16'h73E4: data_out = 8'hF;
                    16'h73E5: data_out = 8'hE;
                    16'h73E6: data_out = 8'hD;
                    16'h73E7: data_out = 8'hC;
                    16'h73E8: data_out = 8'hB;
                    16'h73E9: data_out = 8'hA;
                    16'h73EA: data_out = 8'h9;
                    16'h73EB: data_out = 8'h8;
                    16'h73EC: data_out = 8'h7;
                    16'h73ED: data_out = 8'h6;
                    16'h73EE: data_out = 8'h5;
                    16'h73EF: data_out = 8'h4;
                    16'h73F0: data_out = 8'h3;
                    16'h73F1: data_out = 8'h2;
                    16'h73F2: data_out = 8'h1;
                    16'h73F3: data_out = 8'h0;
                    16'h73F4: data_out = 8'h81;
                    16'h73F5: data_out = 8'h82;
                    16'h73F6: data_out = 8'h83;
                    16'h73F7: data_out = 8'h84;
                    16'h73F8: data_out = 8'h85;
                    16'h73F9: data_out = 8'h86;
                    16'h73FA: data_out = 8'h87;
                    16'h73FB: data_out = 8'h88;
                    16'h73FC: data_out = 8'h89;
                    16'h73FD: data_out = 8'h8A;
                    16'h73FE: data_out = 8'h8B;
                    16'h73FF: data_out = 8'h8C;
                    16'h7400: data_out = 8'h74;
                    16'h7401: data_out = 8'h75;
                    16'h7402: data_out = 8'h76;
                    16'h7403: data_out = 8'h77;
                    16'h7404: data_out = 8'h78;
                    16'h7405: data_out = 8'h79;
                    16'h7406: data_out = 8'h7A;
                    16'h7407: data_out = 8'h7B;
                    16'h7408: data_out = 8'h7C;
                    16'h7409: data_out = 8'h7D;
                    16'h740A: data_out = 8'h7E;
                    16'h740B: data_out = 8'h7F;
                    16'h740C: data_out = 8'h80;
                    16'h740D: data_out = 8'h81;
                    16'h740E: data_out = 8'h82;
                    16'h740F: data_out = 8'h83;
                    16'h7410: data_out = 8'h84;
                    16'h7411: data_out = 8'h85;
                    16'h7412: data_out = 8'h86;
                    16'h7413: data_out = 8'h87;
                    16'h7414: data_out = 8'h88;
                    16'h7415: data_out = 8'h89;
                    16'h7416: data_out = 8'h8A;
                    16'h7417: data_out = 8'h8B;
                    16'h7418: data_out = 8'h8C;
                    16'h7419: data_out = 8'h8D;
                    16'h741A: data_out = 8'h8E;
                    16'h741B: data_out = 8'h8F;
                    16'h741C: data_out = 8'h90;
                    16'h741D: data_out = 8'h91;
                    16'h741E: data_out = 8'h92;
                    16'h741F: data_out = 8'h93;
                    16'h7420: data_out = 8'h94;
                    16'h7421: data_out = 8'h95;
                    16'h7422: data_out = 8'h96;
                    16'h7423: data_out = 8'h97;
                    16'h7424: data_out = 8'h98;
                    16'h7425: data_out = 8'h99;
                    16'h7426: data_out = 8'h9A;
                    16'h7427: data_out = 8'h9B;
                    16'h7428: data_out = 8'h9C;
                    16'h7429: data_out = 8'h9D;
                    16'h742A: data_out = 8'h9E;
                    16'h742B: data_out = 8'h9F;
                    16'h742C: data_out = 8'hA0;
                    16'h742D: data_out = 8'hA1;
                    16'h742E: data_out = 8'hA2;
                    16'h742F: data_out = 8'hA3;
                    16'h7430: data_out = 8'hA4;
                    16'h7431: data_out = 8'hA5;
                    16'h7432: data_out = 8'hA6;
                    16'h7433: data_out = 8'hA7;
                    16'h7434: data_out = 8'hA8;
                    16'h7435: data_out = 8'hA9;
                    16'h7436: data_out = 8'hAA;
                    16'h7437: data_out = 8'hAB;
                    16'h7438: data_out = 8'hAC;
                    16'h7439: data_out = 8'hAD;
                    16'h743A: data_out = 8'hAE;
                    16'h743B: data_out = 8'hAF;
                    16'h743C: data_out = 8'hB0;
                    16'h743D: data_out = 8'hB1;
                    16'h743E: data_out = 8'hB2;
                    16'h743F: data_out = 8'hB3;
                    16'h7440: data_out = 8'hB4;
                    16'h7441: data_out = 8'hB5;
                    16'h7442: data_out = 8'hB6;
                    16'h7443: data_out = 8'hB7;
                    16'h7444: data_out = 8'hB8;
                    16'h7445: data_out = 8'hB9;
                    16'h7446: data_out = 8'hBA;
                    16'h7447: data_out = 8'hBB;
                    16'h7448: data_out = 8'hBC;
                    16'h7449: data_out = 8'hBD;
                    16'h744A: data_out = 8'hBE;
                    16'h744B: data_out = 8'hBF;
                    16'h744C: data_out = 8'hC0;
                    16'h744D: data_out = 8'hC1;
                    16'h744E: data_out = 8'hC2;
                    16'h744F: data_out = 8'hC3;
                    16'h7450: data_out = 8'hC4;
                    16'h7451: data_out = 8'hC5;
                    16'h7452: data_out = 8'hC6;
                    16'h7453: data_out = 8'hC7;
                    16'h7454: data_out = 8'hC8;
                    16'h7455: data_out = 8'hC9;
                    16'h7456: data_out = 8'hCA;
                    16'h7457: data_out = 8'hCB;
                    16'h7458: data_out = 8'hCC;
                    16'h7459: data_out = 8'hCD;
                    16'h745A: data_out = 8'hCE;
                    16'h745B: data_out = 8'hCF;
                    16'h745C: data_out = 8'hD0;
                    16'h745D: data_out = 8'hD1;
                    16'h745E: data_out = 8'hD2;
                    16'h745F: data_out = 8'hD3;
                    16'h7460: data_out = 8'hD4;
                    16'h7461: data_out = 8'hD5;
                    16'h7462: data_out = 8'hD6;
                    16'h7463: data_out = 8'hD7;
                    16'h7464: data_out = 8'hD8;
                    16'h7465: data_out = 8'hD9;
                    16'h7466: data_out = 8'hDA;
                    16'h7467: data_out = 8'hDB;
                    16'h7468: data_out = 8'hDC;
                    16'h7469: data_out = 8'hDD;
                    16'h746A: data_out = 8'hDE;
                    16'h746B: data_out = 8'hDF;
                    16'h746C: data_out = 8'hE0;
                    16'h746D: data_out = 8'hE1;
                    16'h746E: data_out = 8'hE2;
                    16'h746F: data_out = 8'hE3;
                    16'h7470: data_out = 8'hE4;
                    16'h7471: data_out = 8'hE5;
                    16'h7472: data_out = 8'hE6;
                    16'h7473: data_out = 8'hE7;
                    16'h7474: data_out = 8'hE8;
                    16'h7475: data_out = 8'hE9;
                    16'h7476: data_out = 8'hEA;
                    16'h7477: data_out = 8'hEB;
                    16'h7478: data_out = 8'hEC;
                    16'h7479: data_out = 8'hED;
                    16'h747A: data_out = 8'hEE;
                    16'h747B: data_out = 8'hEF;
                    16'h747C: data_out = 8'hF0;
                    16'h747D: data_out = 8'hF1;
                    16'h747E: data_out = 8'hF2;
                    16'h747F: data_out = 8'hF3;
                    16'h7480: data_out = 8'h74;
                    16'h7481: data_out = 8'h73;
                    16'h7482: data_out = 8'h72;
                    16'h7483: data_out = 8'h71;
                    16'h7484: data_out = 8'h70;
                    16'h7485: data_out = 8'h6F;
                    16'h7486: data_out = 8'h6E;
                    16'h7487: data_out = 8'h6D;
                    16'h7488: data_out = 8'h6C;
                    16'h7489: data_out = 8'h6B;
                    16'h748A: data_out = 8'h6A;
                    16'h748B: data_out = 8'h69;
                    16'h748C: data_out = 8'h68;
                    16'h748D: data_out = 8'h67;
                    16'h748E: data_out = 8'h66;
                    16'h748F: data_out = 8'h65;
                    16'h7490: data_out = 8'h64;
                    16'h7491: data_out = 8'h63;
                    16'h7492: data_out = 8'h62;
                    16'h7493: data_out = 8'h61;
                    16'h7494: data_out = 8'h60;
                    16'h7495: data_out = 8'h5F;
                    16'h7496: data_out = 8'h5E;
                    16'h7497: data_out = 8'h5D;
                    16'h7498: data_out = 8'h5C;
                    16'h7499: data_out = 8'h5B;
                    16'h749A: data_out = 8'h5A;
                    16'h749B: data_out = 8'h59;
                    16'h749C: data_out = 8'h58;
                    16'h749D: data_out = 8'h57;
                    16'h749E: data_out = 8'h56;
                    16'h749F: data_out = 8'h55;
                    16'h74A0: data_out = 8'h54;
                    16'h74A1: data_out = 8'h53;
                    16'h74A2: data_out = 8'h52;
                    16'h74A3: data_out = 8'h51;
                    16'h74A4: data_out = 8'h50;
                    16'h74A5: data_out = 8'h4F;
                    16'h74A6: data_out = 8'h4E;
                    16'h74A7: data_out = 8'h4D;
                    16'h74A8: data_out = 8'h4C;
                    16'h74A9: data_out = 8'h4B;
                    16'h74AA: data_out = 8'h4A;
                    16'h74AB: data_out = 8'h49;
                    16'h74AC: data_out = 8'h48;
                    16'h74AD: data_out = 8'h47;
                    16'h74AE: data_out = 8'h46;
                    16'h74AF: data_out = 8'h45;
                    16'h74B0: data_out = 8'h44;
                    16'h74B1: data_out = 8'h43;
                    16'h74B2: data_out = 8'h42;
                    16'h74B3: data_out = 8'h41;
                    16'h74B4: data_out = 8'h40;
                    16'h74B5: data_out = 8'h3F;
                    16'h74B6: data_out = 8'h3E;
                    16'h74B7: data_out = 8'h3D;
                    16'h74B8: data_out = 8'h3C;
                    16'h74B9: data_out = 8'h3B;
                    16'h74BA: data_out = 8'h3A;
                    16'h74BB: data_out = 8'h39;
                    16'h74BC: data_out = 8'h38;
                    16'h74BD: data_out = 8'h37;
                    16'h74BE: data_out = 8'h36;
                    16'h74BF: data_out = 8'h35;
                    16'h74C0: data_out = 8'h34;
                    16'h74C1: data_out = 8'h33;
                    16'h74C2: data_out = 8'h32;
                    16'h74C3: data_out = 8'h31;
                    16'h74C4: data_out = 8'h30;
                    16'h74C5: data_out = 8'h2F;
                    16'h74C6: data_out = 8'h2E;
                    16'h74C7: data_out = 8'h2D;
                    16'h74C8: data_out = 8'h2C;
                    16'h74C9: data_out = 8'h2B;
                    16'h74CA: data_out = 8'h2A;
                    16'h74CB: data_out = 8'h29;
                    16'h74CC: data_out = 8'h28;
                    16'h74CD: data_out = 8'h27;
                    16'h74CE: data_out = 8'h26;
                    16'h74CF: data_out = 8'h25;
                    16'h74D0: data_out = 8'h24;
                    16'h74D1: data_out = 8'h23;
                    16'h74D2: data_out = 8'h22;
                    16'h74D3: data_out = 8'h21;
                    16'h74D4: data_out = 8'h20;
                    16'h74D5: data_out = 8'h1F;
                    16'h74D6: data_out = 8'h1E;
                    16'h74D7: data_out = 8'h1D;
                    16'h74D8: data_out = 8'h1C;
                    16'h74D9: data_out = 8'h1B;
                    16'h74DA: data_out = 8'h1A;
                    16'h74DB: data_out = 8'h19;
                    16'h74DC: data_out = 8'h18;
                    16'h74DD: data_out = 8'h17;
                    16'h74DE: data_out = 8'h16;
                    16'h74DF: data_out = 8'h15;
                    16'h74E0: data_out = 8'h14;
                    16'h74E1: data_out = 8'h13;
                    16'h74E2: data_out = 8'h12;
                    16'h74E3: data_out = 8'h11;
                    16'h74E4: data_out = 8'h10;
                    16'h74E5: data_out = 8'hF;
                    16'h74E6: data_out = 8'hE;
                    16'h74E7: data_out = 8'hD;
                    16'h74E8: data_out = 8'hC;
                    16'h74E9: data_out = 8'hB;
                    16'h74EA: data_out = 8'hA;
                    16'h74EB: data_out = 8'h9;
                    16'h74EC: data_out = 8'h8;
                    16'h74ED: data_out = 8'h7;
                    16'h74EE: data_out = 8'h6;
                    16'h74EF: data_out = 8'h5;
                    16'h74F0: data_out = 8'h4;
                    16'h74F1: data_out = 8'h3;
                    16'h74F2: data_out = 8'h2;
                    16'h74F3: data_out = 8'h1;
                    16'h74F4: data_out = 8'h0;
                    16'h74F5: data_out = 8'h81;
                    16'h74F6: data_out = 8'h82;
                    16'h74F7: data_out = 8'h83;
                    16'h74F8: data_out = 8'h84;
                    16'h74F9: data_out = 8'h85;
                    16'h74FA: data_out = 8'h86;
                    16'h74FB: data_out = 8'h87;
                    16'h74FC: data_out = 8'h88;
                    16'h74FD: data_out = 8'h89;
                    16'h74FE: data_out = 8'h8A;
                    16'h74FF: data_out = 8'h8B;
                    16'h7500: data_out = 8'h75;
                    16'h7501: data_out = 8'h76;
                    16'h7502: data_out = 8'h77;
                    16'h7503: data_out = 8'h78;
                    16'h7504: data_out = 8'h79;
                    16'h7505: data_out = 8'h7A;
                    16'h7506: data_out = 8'h7B;
                    16'h7507: data_out = 8'h7C;
                    16'h7508: data_out = 8'h7D;
                    16'h7509: data_out = 8'h7E;
                    16'h750A: data_out = 8'h7F;
                    16'h750B: data_out = 8'h80;
                    16'h750C: data_out = 8'h81;
                    16'h750D: data_out = 8'h82;
                    16'h750E: data_out = 8'h83;
                    16'h750F: data_out = 8'h84;
                    16'h7510: data_out = 8'h85;
                    16'h7511: data_out = 8'h86;
                    16'h7512: data_out = 8'h87;
                    16'h7513: data_out = 8'h88;
                    16'h7514: data_out = 8'h89;
                    16'h7515: data_out = 8'h8A;
                    16'h7516: data_out = 8'h8B;
                    16'h7517: data_out = 8'h8C;
                    16'h7518: data_out = 8'h8D;
                    16'h7519: data_out = 8'h8E;
                    16'h751A: data_out = 8'h8F;
                    16'h751B: data_out = 8'h90;
                    16'h751C: data_out = 8'h91;
                    16'h751D: data_out = 8'h92;
                    16'h751E: data_out = 8'h93;
                    16'h751F: data_out = 8'h94;
                    16'h7520: data_out = 8'h95;
                    16'h7521: data_out = 8'h96;
                    16'h7522: data_out = 8'h97;
                    16'h7523: data_out = 8'h98;
                    16'h7524: data_out = 8'h99;
                    16'h7525: data_out = 8'h9A;
                    16'h7526: data_out = 8'h9B;
                    16'h7527: data_out = 8'h9C;
                    16'h7528: data_out = 8'h9D;
                    16'h7529: data_out = 8'h9E;
                    16'h752A: data_out = 8'h9F;
                    16'h752B: data_out = 8'hA0;
                    16'h752C: data_out = 8'hA1;
                    16'h752D: data_out = 8'hA2;
                    16'h752E: data_out = 8'hA3;
                    16'h752F: data_out = 8'hA4;
                    16'h7530: data_out = 8'hA5;
                    16'h7531: data_out = 8'hA6;
                    16'h7532: data_out = 8'hA7;
                    16'h7533: data_out = 8'hA8;
                    16'h7534: data_out = 8'hA9;
                    16'h7535: data_out = 8'hAA;
                    16'h7536: data_out = 8'hAB;
                    16'h7537: data_out = 8'hAC;
                    16'h7538: data_out = 8'hAD;
                    16'h7539: data_out = 8'hAE;
                    16'h753A: data_out = 8'hAF;
                    16'h753B: data_out = 8'hB0;
                    16'h753C: data_out = 8'hB1;
                    16'h753D: data_out = 8'hB2;
                    16'h753E: data_out = 8'hB3;
                    16'h753F: data_out = 8'hB4;
                    16'h7540: data_out = 8'hB5;
                    16'h7541: data_out = 8'hB6;
                    16'h7542: data_out = 8'hB7;
                    16'h7543: data_out = 8'hB8;
                    16'h7544: data_out = 8'hB9;
                    16'h7545: data_out = 8'hBA;
                    16'h7546: data_out = 8'hBB;
                    16'h7547: data_out = 8'hBC;
                    16'h7548: data_out = 8'hBD;
                    16'h7549: data_out = 8'hBE;
                    16'h754A: data_out = 8'hBF;
                    16'h754B: data_out = 8'hC0;
                    16'h754C: data_out = 8'hC1;
                    16'h754D: data_out = 8'hC2;
                    16'h754E: data_out = 8'hC3;
                    16'h754F: data_out = 8'hC4;
                    16'h7550: data_out = 8'hC5;
                    16'h7551: data_out = 8'hC6;
                    16'h7552: data_out = 8'hC7;
                    16'h7553: data_out = 8'hC8;
                    16'h7554: data_out = 8'hC9;
                    16'h7555: data_out = 8'hCA;
                    16'h7556: data_out = 8'hCB;
                    16'h7557: data_out = 8'hCC;
                    16'h7558: data_out = 8'hCD;
                    16'h7559: data_out = 8'hCE;
                    16'h755A: data_out = 8'hCF;
                    16'h755B: data_out = 8'hD0;
                    16'h755C: data_out = 8'hD1;
                    16'h755D: data_out = 8'hD2;
                    16'h755E: data_out = 8'hD3;
                    16'h755F: data_out = 8'hD4;
                    16'h7560: data_out = 8'hD5;
                    16'h7561: data_out = 8'hD6;
                    16'h7562: data_out = 8'hD7;
                    16'h7563: data_out = 8'hD8;
                    16'h7564: data_out = 8'hD9;
                    16'h7565: data_out = 8'hDA;
                    16'h7566: data_out = 8'hDB;
                    16'h7567: data_out = 8'hDC;
                    16'h7568: data_out = 8'hDD;
                    16'h7569: data_out = 8'hDE;
                    16'h756A: data_out = 8'hDF;
                    16'h756B: data_out = 8'hE0;
                    16'h756C: data_out = 8'hE1;
                    16'h756D: data_out = 8'hE2;
                    16'h756E: data_out = 8'hE3;
                    16'h756F: data_out = 8'hE4;
                    16'h7570: data_out = 8'hE5;
                    16'h7571: data_out = 8'hE6;
                    16'h7572: data_out = 8'hE7;
                    16'h7573: data_out = 8'hE8;
                    16'h7574: data_out = 8'hE9;
                    16'h7575: data_out = 8'hEA;
                    16'h7576: data_out = 8'hEB;
                    16'h7577: data_out = 8'hEC;
                    16'h7578: data_out = 8'hED;
                    16'h7579: data_out = 8'hEE;
                    16'h757A: data_out = 8'hEF;
                    16'h757B: data_out = 8'hF0;
                    16'h757C: data_out = 8'hF1;
                    16'h757D: data_out = 8'hF2;
                    16'h757E: data_out = 8'hF3;
                    16'h757F: data_out = 8'hF4;
                    16'h7580: data_out = 8'h75;
                    16'h7581: data_out = 8'h74;
                    16'h7582: data_out = 8'h73;
                    16'h7583: data_out = 8'h72;
                    16'h7584: data_out = 8'h71;
                    16'h7585: data_out = 8'h70;
                    16'h7586: data_out = 8'h6F;
                    16'h7587: data_out = 8'h6E;
                    16'h7588: data_out = 8'h6D;
                    16'h7589: data_out = 8'h6C;
                    16'h758A: data_out = 8'h6B;
                    16'h758B: data_out = 8'h6A;
                    16'h758C: data_out = 8'h69;
                    16'h758D: data_out = 8'h68;
                    16'h758E: data_out = 8'h67;
                    16'h758F: data_out = 8'h66;
                    16'h7590: data_out = 8'h65;
                    16'h7591: data_out = 8'h64;
                    16'h7592: data_out = 8'h63;
                    16'h7593: data_out = 8'h62;
                    16'h7594: data_out = 8'h61;
                    16'h7595: data_out = 8'h60;
                    16'h7596: data_out = 8'h5F;
                    16'h7597: data_out = 8'h5E;
                    16'h7598: data_out = 8'h5D;
                    16'h7599: data_out = 8'h5C;
                    16'h759A: data_out = 8'h5B;
                    16'h759B: data_out = 8'h5A;
                    16'h759C: data_out = 8'h59;
                    16'h759D: data_out = 8'h58;
                    16'h759E: data_out = 8'h57;
                    16'h759F: data_out = 8'h56;
                    16'h75A0: data_out = 8'h55;
                    16'h75A1: data_out = 8'h54;
                    16'h75A2: data_out = 8'h53;
                    16'h75A3: data_out = 8'h52;
                    16'h75A4: data_out = 8'h51;
                    16'h75A5: data_out = 8'h50;
                    16'h75A6: data_out = 8'h4F;
                    16'h75A7: data_out = 8'h4E;
                    16'h75A8: data_out = 8'h4D;
                    16'h75A9: data_out = 8'h4C;
                    16'h75AA: data_out = 8'h4B;
                    16'h75AB: data_out = 8'h4A;
                    16'h75AC: data_out = 8'h49;
                    16'h75AD: data_out = 8'h48;
                    16'h75AE: data_out = 8'h47;
                    16'h75AF: data_out = 8'h46;
                    16'h75B0: data_out = 8'h45;
                    16'h75B1: data_out = 8'h44;
                    16'h75B2: data_out = 8'h43;
                    16'h75B3: data_out = 8'h42;
                    16'h75B4: data_out = 8'h41;
                    16'h75B5: data_out = 8'h40;
                    16'h75B6: data_out = 8'h3F;
                    16'h75B7: data_out = 8'h3E;
                    16'h75B8: data_out = 8'h3D;
                    16'h75B9: data_out = 8'h3C;
                    16'h75BA: data_out = 8'h3B;
                    16'h75BB: data_out = 8'h3A;
                    16'h75BC: data_out = 8'h39;
                    16'h75BD: data_out = 8'h38;
                    16'h75BE: data_out = 8'h37;
                    16'h75BF: data_out = 8'h36;
                    16'h75C0: data_out = 8'h35;
                    16'h75C1: data_out = 8'h34;
                    16'h75C2: data_out = 8'h33;
                    16'h75C3: data_out = 8'h32;
                    16'h75C4: data_out = 8'h31;
                    16'h75C5: data_out = 8'h30;
                    16'h75C6: data_out = 8'h2F;
                    16'h75C7: data_out = 8'h2E;
                    16'h75C8: data_out = 8'h2D;
                    16'h75C9: data_out = 8'h2C;
                    16'h75CA: data_out = 8'h2B;
                    16'h75CB: data_out = 8'h2A;
                    16'h75CC: data_out = 8'h29;
                    16'h75CD: data_out = 8'h28;
                    16'h75CE: data_out = 8'h27;
                    16'h75CF: data_out = 8'h26;
                    16'h75D0: data_out = 8'h25;
                    16'h75D1: data_out = 8'h24;
                    16'h75D2: data_out = 8'h23;
                    16'h75D3: data_out = 8'h22;
                    16'h75D4: data_out = 8'h21;
                    16'h75D5: data_out = 8'h20;
                    16'h75D6: data_out = 8'h1F;
                    16'h75D7: data_out = 8'h1E;
                    16'h75D8: data_out = 8'h1D;
                    16'h75D9: data_out = 8'h1C;
                    16'h75DA: data_out = 8'h1B;
                    16'h75DB: data_out = 8'h1A;
                    16'h75DC: data_out = 8'h19;
                    16'h75DD: data_out = 8'h18;
                    16'h75DE: data_out = 8'h17;
                    16'h75DF: data_out = 8'h16;
                    16'h75E0: data_out = 8'h15;
                    16'h75E1: data_out = 8'h14;
                    16'h75E2: data_out = 8'h13;
                    16'h75E3: data_out = 8'h12;
                    16'h75E4: data_out = 8'h11;
                    16'h75E5: data_out = 8'h10;
                    16'h75E6: data_out = 8'hF;
                    16'h75E7: data_out = 8'hE;
                    16'h75E8: data_out = 8'hD;
                    16'h75E9: data_out = 8'hC;
                    16'h75EA: data_out = 8'hB;
                    16'h75EB: data_out = 8'hA;
                    16'h75EC: data_out = 8'h9;
                    16'h75ED: data_out = 8'h8;
                    16'h75EE: data_out = 8'h7;
                    16'h75EF: data_out = 8'h6;
                    16'h75F0: data_out = 8'h5;
                    16'h75F1: data_out = 8'h4;
                    16'h75F2: data_out = 8'h3;
                    16'h75F3: data_out = 8'h2;
                    16'h75F4: data_out = 8'h1;
                    16'h75F5: data_out = 8'h0;
                    16'h75F6: data_out = 8'h81;
                    16'h75F7: data_out = 8'h82;
                    16'h75F8: data_out = 8'h83;
                    16'h75F9: data_out = 8'h84;
                    16'h75FA: data_out = 8'h85;
                    16'h75FB: data_out = 8'h86;
                    16'h75FC: data_out = 8'h87;
                    16'h75FD: data_out = 8'h88;
                    16'h75FE: data_out = 8'h89;
                    16'h75FF: data_out = 8'h8A;
                    16'h7600: data_out = 8'h76;
                    16'h7601: data_out = 8'h77;
                    16'h7602: data_out = 8'h78;
                    16'h7603: data_out = 8'h79;
                    16'h7604: data_out = 8'h7A;
                    16'h7605: data_out = 8'h7B;
                    16'h7606: data_out = 8'h7C;
                    16'h7607: data_out = 8'h7D;
                    16'h7608: data_out = 8'h7E;
                    16'h7609: data_out = 8'h7F;
                    16'h760A: data_out = 8'h80;
                    16'h760B: data_out = 8'h81;
                    16'h760C: data_out = 8'h82;
                    16'h760D: data_out = 8'h83;
                    16'h760E: data_out = 8'h84;
                    16'h760F: data_out = 8'h85;
                    16'h7610: data_out = 8'h86;
                    16'h7611: data_out = 8'h87;
                    16'h7612: data_out = 8'h88;
                    16'h7613: data_out = 8'h89;
                    16'h7614: data_out = 8'h8A;
                    16'h7615: data_out = 8'h8B;
                    16'h7616: data_out = 8'h8C;
                    16'h7617: data_out = 8'h8D;
                    16'h7618: data_out = 8'h8E;
                    16'h7619: data_out = 8'h8F;
                    16'h761A: data_out = 8'h90;
                    16'h761B: data_out = 8'h91;
                    16'h761C: data_out = 8'h92;
                    16'h761D: data_out = 8'h93;
                    16'h761E: data_out = 8'h94;
                    16'h761F: data_out = 8'h95;
                    16'h7620: data_out = 8'h96;
                    16'h7621: data_out = 8'h97;
                    16'h7622: data_out = 8'h98;
                    16'h7623: data_out = 8'h99;
                    16'h7624: data_out = 8'h9A;
                    16'h7625: data_out = 8'h9B;
                    16'h7626: data_out = 8'h9C;
                    16'h7627: data_out = 8'h9D;
                    16'h7628: data_out = 8'h9E;
                    16'h7629: data_out = 8'h9F;
                    16'h762A: data_out = 8'hA0;
                    16'h762B: data_out = 8'hA1;
                    16'h762C: data_out = 8'hA2;
                    16'h762D: data_out = 8'hA3;
                    16'h762E: data_out = 8'hA4;
                    16'h762F: data_out = 8'hA5;
                    16'h7630: data_out = 8'hA6;
                    16'h7631: data_out = 8'hA7;
                    16'h7632: data_out = 8'hA8;
                    16'h7633: data_out = 8'hA9;
                    16'h7634: data_out = 8'hAA;
                    16'h7635: data_out = 8'hAB;
                    16'h7636: data_out = 8'hAC;
                    16'h7637: data_out = 8'hAD;
                    16'h7638: data_out = 8'hAE;
                    16'h7639: data_out = 8'hAF;
                    16'h763A: data_out = 8'hB0;
                    16'h763B: data_out = 8'hB1;
                    16'h763C: data_out = 8'hB2;
                    16'h763D: data_out = 8'hB3;
                    16'h763E: data_out = 8'hB4;
                    16'h763F: data_out = 8'hB5;
                    16'h7640: data_out = 8'hB6;
                    16'h7641: data_out = 8'hB7;
                    16'h7642: data_out = 8'hB8;
                    16'h7643: data_out = 8'hB9;
                    16'h7644: data_out = 8'hBA;
                    16'h7645: data_out = 8'hBB;
                    16'h7646: data_out = 8'hBC;
                    16'h7647: data_out = 8'hBD;
                    16'h7648: data_out = 8'hBE;
                    16'h7649: data_out = 8'hBF;
                    16'h764A: data_out = 8'hC0;
                    16'h764B: data_out = 8'hC1;
                    16'h764C: data_out = 8'hC2;
                    16'h764D: data_out = 8'hC3;
                    16'h764E: data_out = 8'hC4;
                    16'h764F: data_out = 8'hC5;
                    16'h7650: data_out = 8'hC6;
                    16'h7651: data_out = 8'hC7;
                    16'h7652: data_out = 8'hC8;
                    16'h7653: data_out = 8'hC9;
                    16'h7654: data_out = 8'hCA;
                    16'h7655: data_out = 8'hCB;
                    16'h7656: data_out = 8'hCC;
                    16'h7657: data_out = 8'hCD;
                    16'h7658: data_out = 8'hCE;
                    16'h7659: data_out = 8'hCF;
                    16'h765A: data_out = 8'hD0;
                    16'h765B: data_out = 8'hD1;
                    16'h765C: data_out = 8'hD2;
                    16'h765D: data_out = 8'hD3;
                    16'h765E: data_out = 8'hD4;
                    16'h765F: data_out = 8'hD5;
                    16'h7660: data_out = 8'hD6;
                    16'h7661: data_out = 8'hD7;
                    16'h7662: data_out = 8'hD8;
                    16'h7663: data_out = 8'hD9;
                    16'h7664: data_out = 8'hDA;
                    16'h7665: data_out = 8'hDB;
                    16'h7666: data_out = 8'hDC;
                    16'h7667: data_out = 8'hDD;
                    16'h7668: data_out = 8'hDE;
                    16'h7669: data_out = 8'hDF;
                    16'h766A: data_out = 8'hE0;
                    16'h766B: data_out = 8'hE1;
                    16'h766C: data_out = 8'hE2;
                    16'h766D: data_out = 8'hE3;
                    16'h766E: data_out = 8'hE4;
                    16'h766F: data_out = 8'hE5;
                    16'h7670: data_out = 8'hE6;
                    16'h7671: data_out = 8'hE7;
                    16'h7672: data_out = 8'hE8;
                    16'h7673: data_out = 8'hE9;
                    16'h7674: data_out = 8'hEA;
                    16'h7675: data_out = 8'hEB;
                    16'h7676: data_out = 8'hEC;
                    16'h7677: data_out = 8'hED;
                    16'h7678: data_out = 8'hEE;
                    16'h7679: data_out = 8'hEF;
                    16'h767A: data_out = 8'hF0;
                    16'h767B: data_out = 8'hF1;
                    16'h767C: data_out = 8'hF2;
                    16'h767D: data_out = 8'hF3;
                    16'h767E: data_out = 8'hF4;
                    16'h767F: data_out = 8'hF5;
                    16'h7680: data_out = 8'h76;
                    16'h7681: data_out = 8'h75;
                    16'h7682: data_out = 8'h74;
                    16'h7683: data_out = 8'h73;
                    16'h7684: data_out = 8'h72;
                    16'h7685: data_out = 8'h71;
                    16'h7686: data_out = 8'h70;
                    16'h7687: data_out = 8'h6F;
                    16'h7688: data_out = 8'h6E;
                    16'h7689: data_out = 8'h6D;
                    16'h768A: data_out = 8'h6C;
                    16'h768B: data_out = 8'h6B;
                    16'h768C: data_out = 8'h6A;
                    16'h768D: data_out = 8'h69;
                    16'h768E: data_out = 8'h68;
                    16'h768F: data_out = 8'h67;
                    16'h7690: data_out = 8'h66;
                    16'h7691: data_out = 8'h65;
                    16'h7692: data_out = 8'h64;
                    16'h7693: data_out = 8'h63;
                    16'h7694: data_out = 8'h62;
                    16'h7695: data_out = 8'h61;
                    16'h7696: data_out = 8'h60;
                    16'h7697: data_out = 8'h5F;
                    16'h7698: data_out = 8'h5E;
                    16'h7699: data_out = 8'h5D;
                    16'h769A: data_out = 8'h5C;
                    16'h769B: data_out = 8'h5B;
                    16'h769C: data_out = 8'h5A;
                    16'h769D: data_out = 8'h59;
                    16'h769E: data_out = 8'h58;
                    16'h769F: data_out = 8'h57;
                    16'h76A0: data_out = 8'h56;
                    16'h76A1: data_out = 8'h55;
                    16'h76A2: data_out = 8'h54;
                    16'h76A3: data_out = 8'h53;
                    16'h76A4: data_out = 8'h52;
                    16'h76A5: data_out = 8'h51;
                    16'h76A6: data_out = 8'h50;
                    16'h76A7: data_out = 8'h4F;
                    16'h76A8: data_out = 8'h4E;
                    16'h76A9: data_out = 8'h4D;
                    16'h76AA: data_out = 8'h4C;
                    16'h76AB: data_out = 8'h4B;
                    16'h76AC: data_out = 8'h4A;
                    16'h76AD: data_out = 8'h49;
                    16'h76AE: data_out = 8'h48;
                    16'h76AF: data_out = 8'h47;
                    16'h76B0: data_out = 8'h46;
                    16'h76B1: data_out = 8'h45;
                    16'h76B2: data_out = 8'h44;
                    16'h76B3: data_out = 8'h43;
                    16'h76B4: data_out = 8'h42;
                    16'h76B5: data_out = 8'h41;
                    16'h76B6: data_out = 8'h40;
                    16'h76B7: data_out = 8'h3F;
                    16'h76B8: data_out = 8'h3E;
                    16'h76B9: data_out = 8'h3D;
                    16'h76BA: data_out = 8'h3C;
                    16'h76BB: data_out = 8'h3B;
                    16'h76BC: data_out = 8'h3A;
                    16'h76BD: data_out = 8'h39;
                    16'h76BE: data_out = 8'h38;
                    16'h76BF: data_out = 8'h37;
                    16'h76C0: data_out = 8'h36;
                    16'h76C1: data_out = 8'h35;
                    16'h76C2: data_out = 8'h34;
                    16'h76C3: data_out = 8'h33;
                    16'h76C4: data_out = 8'h32;
                    16'h76C5: data_out = 8'h31;
                    16'h76C6: data_out = 8'h30;
                    16'h76C7: data_out = 8'h2F;
                    16'h76C8: data_out = 8'h2E;
                    16'h76C9: data_out = 8'h2D;
                    16'h76CA: data_out = 8'h2C;
                    16'h76CB: data_out = 8'h2B;
                    16'h76CC: data_out = 8'h2A;
                    16'h76CD: data_out = 8'h29;
                    16'h76CE: data_out = 8'h28;
                    16'h76CF: data_out = 8'h27;
                    16'h76D0: data_out = 8'h26;
                    16'h76D1: data_out = 8'h25;
                    16'h76D2: data_out = 8'h24;
                    16'h76D3: data_out = 8'h23;
                    16'h76D4: data_out = 8'h22;
                    16'h76D5: data_out = 8'h21;
                    16'h76D6: data_out = 8'h20;
                    16'h76D7: data_out = 8'h1F;
                    16'h76D8: data_out = 8'h1E;
                    16'h76D9: data_out = 8'h1D;
                    16'h76DA: data_out = 8'h1C;
                    16'h76DB: data_out = 8'h1B;
                    16'h76DC: data_out = 8'h1A;
                    16'h76DD: data_out = 8'h19;
                    16'h76DE: data_out = 8'h18;
                    16'h76DF: data_out = 8'h17;
                    16'h76E0: data_out = 8'h16;
                    16'h76E1: data_out = 8'h15;
                    16'h76E2: data_out = 8'h14;
                    16'h76E3: data_out = 8'h13;
                    16'h76E4: data_out = 8'h12;
                    16'h76E5: data_out = 8'h11;
                    16'h76E6: data_out = 8'h10;
                    16'h76E7: data_out = 8'hF;
                    16'h76E8: data_out = 8'hE;
                    16'h76E9: data_out = 8'hD;
                    16'h76EA: data_out = 8'hC;
                    16'h76EB: data_out = 8'hB;
                    16'h76EC: data_out = 8'hA;
                    16'h76ED: data_out = 8'h9;
                    16'h76EE: data_out = 8'h8;
                    16'h76EF: data_out = 8'h7;
                    16'h76F0: data_out = 8'h6;
                    16'h76F1: data_out = 8'h5;
                    16'h76F2: data_out = 8'h4;
                    16'h76F3: data_out = 8'h3;
                    16'h76F4: data_out = 8'h2;
                    16'h76F5: data_out = 8'h1;
                    16'h76F6: data_out = 8'h0;
                    16'h76F7: data_out = 8'h81;
                    16'h76F8: data_out = 8'h82;
                    16'h76F9: data_out = 8'h83;
                    16'h76FA: data_out = 8'h84;
                    16'h76FB: data_out = 8'h85;
                    16'h76FC: data_out = 8'h86;
                    16'h76FD: data_out = 8'h87;
                    16'h76FE: data_out = 8'h88;
                    16'h76FF: data_out = 8'h89;
                    16'h7700: data_out = 8'h77;
                    16'h7701: data_out = 8'h78;
                    16'h7702: data_out = 8'h79;
                    16'h7703: data_out = 8'h7A;
                    16'h7704: data_out = 8'h7B;
                    16'h7705: data_out = 8'h7C;
                    16'h7706: data_out = 8'h7D;
                    16'h7707: data_out = 8'h7E;
                    16'h7708: data_out = 8'h7F;
                    16'h7709: data_out = 8'h80;
                    16'h770A: data_out = 8'h81;
                    16'h770B: data_out = 8'h82;
                    16'h770C: data_out = 8'h83;
                    16'h770D: data_out = 8'h84;
                    16'h770E: data_out = 8'h85;
                    16'h770F: data_out = 8'h86;
                    16'h7710: data_out = 8'h87;
                    16'h7711: data_out = 8'h88;
                    16'h7712: data_out = 8'h89;
                    16'h7713: data_out = 8'h8A;
                    16'h7714: data_out = 8'h8B;
                    16'h7715: data_out = 8'h8C;
                    16'h7716: data_out = 8'h8D;
                    16'h7717: data_out = 8'h8E;
                    16'h7718: data_out = 8'h8F;
                    16'h7719: data_out = 8'h90;
                    16'h771A: data_out = 8'h91;
                    16'h771B: data_out = 8'h92;
                    16'h771C: data_out = 8'h93;
                    16'h771D: data_out = 8'h94;
                    16'h771E: data_out = 8'h95;
                    16'h771F: data_out = 8'h96;
                    16'h7720: data_out = 8'h97;
                    16'h7721: data_out = 8'h98;
                    16'h7722: data_out = 8'h99;
                    16'h7723: data_out = 8'h9A;
                    16'h7724: data_out = 8'h9B;
                    16'h7725: data_out = 8'h9C;
                    16'h7726: data_out = 8'h9D;
                    16'h7727: data_out = 8'h9E;
                    16'h7728: data_out = 8'h9F;
                    16'h7729: data_out = 8'hA0;
                    16'h772A: data_out = 8'hA1;
                    16'h772B: data_out = 8'hA2;
                    16'h772C: data_out = 8'hA3;
                    16'h772D: data_out = 8'hA4;
                    16'h772E: data_out = 8'hA5;
                    16'h772F: data_out = 8'hA6;
                    16'h7730: data_out = 8'hA7;
                    16'h7731: data_out = 8'hA8;
                    16'h7732: data_out = 8'hA9;
                    16'h7733: data_out = 8'hAA;
                    16'h7734: data_out = 8'hAB;
                    16'h7735: data_out = 8'hAC;
                    16'h7736: data_out = 8'hAD;
                    16'h7737: data_out = 8'hAE;
                    16'h7738: data_out = 8'hAF;
                    16'h7739: data_out = 8'hB0;
                    16'h773A: data_out = 8'hB1;
                    16'h773B: data_out = 8'hB2;
                    16'h773C: data_out = 8'hB3;
                    16'h773D: data_out = 8'hB4;
                    16'h773E: data_out = 8'hB5;
                    16'h773F: data_out = 8'hB6;
                    16'h7740: data_out = 8'hB7;
                    16'h7741: data_out = 8'hB8;
                    16'h7742: data_out = 8'hB9;
                    16'h7743: data_out = 8'hBA;
                    16'h7744: data_out = 8'hBB;
                    16'h7745: data_out = 8'hBC;
                    16'h7746: data_out = 8'hBD;
                    16'h7747: data_out = 8'hBE;
                    16'h7748: data_out = 8'hBF;
                    16'h7749: data_out = 8'hC0;
                    16'h774A: data_out = 8'hC1;
                    16'h774B: data_out = 8'hC2;
                    16'h774C: data_out = 8'hC3;
                    16'h774D: data_out = 8'hC4;
                    16'h774E: data_out = 8'hC5;
                    16'h774F: data_out = 8'hC6;
                    16'h7750: data_out = 8'hC7;
                    16'h7751: data_out = 8'hC8;
                    16'h7752: data_out = 8'hC9;
                    16'h7753: data_out = 8'hCA;
                    16'h7754: data_out = 8'hCB;
                    16'h7755: data_out = 8'hCC;
                    16'h7756: data_out = 8'hCD;
                    16'h7757: data_out = 8'hCE;
                    16'h7758: data_out = 8'hCF;
                    16'h7759: data_out = 8'hD0;
                    16'h775A: data_out = 8'hD1;
                    16'h775B: data_out = 8'hD2;
                    16'h775C: data_out = 8'hD3;
                    16'h775D: data_out = 8'hD4;
                    16'h775E: data_out = 8'hD5;
                    16'h775F: data_out = 8'hD6;
                    16'h7760: data_out = 8'hD7;
                    16'h7761: data_out = 8'hD8;
                    16'h7762: data_out = 8'hD9;
                    16'h7763: data_out = 8'hDA;
                    16'h7764: data_out = 8'hDB;
                    16'h7765: data_out = 8'hDC;
                    16'h7766: data_out = 8'hDD;
                    16'h7767: data_out = 8'hDE;
                    16'h7768: data_out = 8'hDF;
                    16'h7769: data_out = 8'hE0;
                    16'h776A: data_out = 8'hE1;
                    16'h776B: data_out = 8'hE2;
                    16'h776C: data_out = 8'hE3;
                    16'h776D: data_out = 8'hE4;
                    16'h776E: data_out = 8'hE5;
                    16'h776F: data_out = 8'hE6;
                    16'h7770: data_out = 8'hE7;
                    16'h7771: data_out = 8'hE8;
                    16'h7772: data_out = 8'hE9;
                    16'h7773: data_out = 8'hEA;
                    16'h7774: data_out = 8'hEB;
                    16'h7775: data_out = 8'hEC;
                    16'h7776: data_out = 8'hED;
                    16'h7777: data_out = 8'hEE;
                    16'h7778: data_out = 8'hEF;
                    16'h7779: data_out = 8'hF0;
                    16'h777A: data_out = 8'hF1;
                    16'h777B: data_out = 8'hF2;
                    16'h777C: data_out = 8'hF3;
                    16'h777D: data_out = 8'hF4;
                    16'h777E: data_out = 8'hF5;
                    16'h777F: data_out = 8'hF6;
                    16'h7780: data_out = 8'h77;
                    16'h7781: data_out = 8'h76;
                    16'h7782: data_out = 8'h75;
                    16'h7783: data_out = 8'h74;
                    16'h7784: data_out = 8'h73;
                    16'h7785: data_out = 8'h72;
                    16'h7786: data_out = 8'h71;
                    16'h7787: data_out = 8'h70;
                    16'h7788: data_out = 8'h6F;
                    16'h7789: data_out = 8'h6E;
                    16'h778A: data_out = 8'h6D;
                    16'h778B: data_out = 8'h6C;
                    16'h778C: data_out = 8'h6B;
                    16'h778D: data_out = 8'h6A;
                    16'h778E: data_out = 8'h69;
                    16'h778F: data_out = 8'h68;
                    16'h7790: data_out = 8'h67;
                    16'h7791: data_out = 8'h66;
                    16'h7792: data_out = 8'h65;
                    16'h7793: data_out = 8'h64;
                    16'h7794: data_out = 8'h63;
                    16'h7795: data_out = 8'h62;
                    16'h7796: data_out = 8'h61;
                    16'h7797: data_out = 8'h60;
                    16'h7798: data_out = 8'h5F;
                    16'h7799: data_out = 8'h5E;
                    16'h779A: data_out = 8'h5D;
                    16'h779B: data_out = 8'h5C;
                    16'h779C: data_out = 8'h5B;
                    16'h779D: data_out = 8'h5A;
                    16'h779E: data_out = 8'h59;
                    16'h779F: data_out = 8'h58;
                    16'h77A0: data_out = 8'h57;
                    16'h77A1: data_out = 8'h56;
                    16'h77A2: data_out = 8'h55;
                    16'h77A3: data_out = 8'h54;
                    16'h77A4: data_out = 8'h53;
                    16'h77A5: data_out = 8'h52;
                    16'h77A6: data_out = 8'h51;
                    16'h77A7: data_out = 8'h50;
                    16'h77A8: data_out = 8'h4F;
                    16'h77A9: data_out = 8'h4E;
                    16'h77AA: data_out = 8'h4D;
                    16'h77AB: data_out = 8'h4C;
                    16'h77AC: data_out = 8'h4B;
                    16'h77AD: data_out = 8'h4A;
                    16'h77AE: data_out = 8'h49;
                    16'h77AF: data_out = 8'h48;
                    16'h77B0: data_out = 8'h47;
                    16'h77B1: data_out = 8'h46;
                    16'h77B2: data_out = 8'h45;
                    16'h77B3: data_out = 8'h44;
                    16'h77B4: data_out = 8'h43;
                    16'h77B5: data_out = 8'h42;
                    16'h77B6: data_out = 8'h41;
                    16'h77B7: data_out = 8'h40;
                    16'h77B8: data_out = 8'h3F;
                    16'h77B9: data_out = 8'h3E;
                    16'h77BA: data_out = 8'h3D;
                    16'h77BB: data_out = 8'h3C;
                    16'h77BC: data_out = 8'h3B;
                    16'h77BD: data_out = 8'h3A;
                    16'h77BE: data_out = 8'h39;
                    16'h77BF: data_out = 8'h38;
                    16'h77C0: data_out = 8'h37;
                    16'h77C1: data_out = 8'h36;
                    16'h77C2: data_out = 8'h35;
                    16'h77C3: data_out = 8'h34;
                    16'h77C4: data_out = 8'h33;
                    16'h77C5: data_out = 8'h32;
                    16'h77C6: data_out = 8'h31;
                    16'h77C7: data_out = 8'h30;
                    16'h77C8: data_out = 8'h2F;
                    16'h77C9: data_out = 8'h2E;
                    16'h77CA: data_out = 8'h2D;
                    16'h77CB: data_out = 8'h2C;
                    16'h77CC: data_out = 8'h2B;
                    16'h77CD: data_out = 8'h2A;
                    16'h77CE: data_out = 8'h29;
                    16'h77CF: data_out = 8'h28;
                    16'h77D0: data_out = 8'h27;
                    16'h77D1: data_out = 8'h26;
                    16'h77D2: data_out = 8'h25;
                    16'h77D3: data_out = 8'h24;
                    16'h77D4: data_out = 8'h23;
                    16'h77D5: data_out = 8'h22;
                    16'h77D6: data_out = 8'h21;
                    16'h77D7: data_out = 8'h20;
                    16'h77D8: data_out = 8'h1F;
                    16'h77D9: data_out = 8'h1E;
                    16'h77DA: data_out = 8'h1D;
                    16'h77DB: data_out = 8'h1C;
                    16'h77DC: data_out = 8'h1B;
                    16'h77DD: data_out = 8'h1A;
                    16'h77DE: data_out = 8'h19;
                    16'h77DF: data_out = 8'h18;
                    16'h77E0: data_out = 8'h17;
                    16'h77E1: data_out = 8'h16;
                    16'h77E2: data_out = 8'h15;
                    16'h77E3: data_out = 8'h14;
                    16'h77E4: data_out = 8'h13;
                    16'h77E5: data_out = 8'h12;
                    16'h77E6: data_out = 8'h11;
                    16'h77E7: data_out = 8'h10;
                    16'h77E8: data_out = 8'hF;
                    16'h77E9: data_out = 8'hE;
                    16'h77EA: data_out = 8'hD;
                    16'h77EB: data_out = 8'hC;
                    16'h77EC: data_out = 8'hB;
                    16'h77ED: data_out = 8'hA;
                    16'h77EE: data_out = 8'h9;
                    16'h77EF: data_out = 8'h8;
                    16'h77F0: data_out = 8'h7;
                    16'h77F1: data_out = 8'h6;
                    16'h77F2: data_out = 8'h5;
                    16'h77F3: data_out = 8'h4;
                    16'h77F4: data_out = 8'h3;
                    16'h77F5: data_out = 8'h2;
                    16'h77F6: data_out = 8'h1;
                    16'h77F7: data_out = 8'h0;
                    16'h77F8: data_out = 8'h81;
                    16'h77F9: data_out = 8'h82;
                    16'h77FA: data_out = 8'h83;
                    16'h77FB: data_out = 8'h84;
                    16'h77FC: data_out = 8'h85;
                    16'h77FD: data_out = 8'h86;
                    16'h77FE: data_out = 8'h87;
                    16'h77FF: data_out = 8'h88;
                    16'h7800: data_out = 8'h78;
                    16'h7801: data_out = 8'h79;
                    16'h7802: data_out = 8'h7A;
                    16'h7803: data_out = 8'h7B;
                    16'h7804: data_out = 8'h7C;
                    16'h7805: data_out = 8'h7D;
                    16'h7806: data_out = 8'h7E;
                    16'h7807: data_out = 8'h7F;
                    16'h7808: data_out = 8'h80;
                    16'h7809: data_out = 8'h81;
                    16'h780A: data_out = 8'h82;
                    16'h780B: data_out = 8'h83;
                    16'h780C: data_out = 8'h84;
                    16'h780D: data_out = 8'h85;
                    16'h780E: data_out = 8'h86;
                    16'h780F: data_out = 8'h87;
                    16'h7810: data_out = 8'h88;
                    16'h7811: data_out = 8'h89;
                    16'h7812: data_out = 8'h8A;
                    16'h7813: data_out = 8'h8B;
                    16'h7814: data_out = 8'h8C;
                    16'h7815: data_out = 8'h8D;
                    16'h7816: data_out = 8'h8E;
                    16'h7817: data_out = 8'h8F;
                    16'h7818: data_out = 8'h90;
                    16'h7819: data_out = 8'h91;
                    16'h781A: data_out = 8'h92;
                    16'h781B: data_out = 8'h93;
                    16'h781C: data_out = 8'h94;
                    16'h781D: data_out = 8'h95;
                    16'h781E: data_out = 8'h96;
                    16'h781F: data_out = 8'h97;
                    16'h7820: data_out = 8'h98;
                    16'h7821: data_out = 8'h99;
                    16'h7822: data_out = 8'h9A;
                    16'h7823: data_out = 8'h9B;
                    16'h7824: data_out = 8'h9C;
                    16'h7825: data_out = 8'h9D;
                    16'h7826: data_out = 8'h9E;
                    16'h7827: data_out = 8'h9F;
                    16'h7828: data_out = 8'hA0;
                    16'h7829: data_out = 8'hA1;
                    16'h782A: data_out = 8'hA2;
                    16'h782B: data_out = 8'hA3;
                    16'h782C: data_out = 8'hA4;
                    16'h782D: data_out = 8'hA5;
                    16'h782E: data_out = 8'hA6;
                    16'h782F: data_out = 8'hA7;
                    16'h7830: data_out = 8'hA8;
                    16'h7831: data_out = 8'hA9;
                    16'h7832: data_out = 8'hAA;
                    16'h7833: data_out = 8'hAB;
                    16'h7834: data_out = 8'hAC;
                    16'h7835: data_out = 8'hAD;
                    16'h7836: data_out = 8'hAE;
                    16'h7837: data_out = 8'hAF;
                    16'h7838: data_out = 8'hB0;
                    16'h7839: data_out = 8'hB1;
                    16'h783A: data_out = 8'hB2;
                    16'h783B: data_out = 8'hB3;
                    16'h783C: data_out = 8'hB4;
                    16'h783D: data_out = 8'hB5;
                    16'h783E: data_out = 8'hB6;
                    16'h783F: data_out = 8'hB7;
                    16'h7840: data_out = 8'hB8;
                    16'h7841: data_out = 8'hB9;
                    16'h7842: data_out = 8'hBA;
                    16'h7843: data_out = 8'hBB;
                    16'h7844: data_out = 8'hBC;
                    16'h7845: data_out = 8'hBD;
                    16'h7846: data_out = 8'hBE;
                    16'h7847: data_out = 8'hBF;
                    16'h7848: data_out = 8'hC0;
                    16'h7849: data_out = 8'hC1;
                    16'h784A: data_out = 8'hC2;
                    16'h784B: data_out = 8'hC3;
                    16'h784C: data_out = 8'hC4;
                    16'h784D: data_out = 8'hC5;
                    16'h784E: data_out = 8'hC6;
                    16'h784F: data_out = 8'hC7;
                    16'h7850: data_out = 8'hC8;
                    16'h7851: data_out = 8'hC9;
                    16'h7852: data_out = 8'hCA;
                    16'h7853: data_out = 8'hCB;
                    16'h7854: data_out = 8'hCC;
                    16'h7855: data_out = 8'hCD;
                    16'h7856: data_out = 8'hCE;
                    16'h7857: data_out = 8'hCF;
                    16'h7858: data_out = 8'hD0;
                    16'h7859: data_out = 8'hD1;
                    16'h785A: data_out = 8'hD2;
                    16'h785B: data_out = 8'hD3;
                    16'h785C: data_out = 8'hD4;
                    16'h785D: data_out = 8'hD5;
                    16'h785E: data_out = 8'hD6;
                    16'h785F: data_out = 8'hD7;
                    16'h7860: data_out = 8'hD8;
                    16'h7861: data_out = 8'hD9;
                    16'h7862: data_out = 8'hDA;
                    16'h7863: data_out = 8'hDB;
                    16'h7864: data_out = 8'hDC;
                    16'h7865: data_out = 8'hDD;
                    16'h7866: data_out = 8'hDE;
                    16'h7867: data_out = 8'hDF;
                    16'h7868: data_out = 8'hE0;
                    16'h7869: data_out = 8'hE1;
                    16'h786A: data_out = 8'hE2;
                    16'h786B: data_out = 8'hE3;
                    16'h786C: data_out = 8'hE4;
                    16'h786D: data_out = 8'hE5;
                    16'h786E: data_out = 8'hE6;
                    16'h786F: data_out = 8'hE7;
                    16'h7870: data_out = 8'hE8;
                    16'h7871: data_out = 8'hE9;
                    16'h7872: data_out = 8'hEA;
                    16'h7873: data_out = 8'hEB;
                    16'h7874: data_out = 8'hEC;
                    16'h7875: data_out = 8'hED;
                    16'h7876: data_out = 8'hEE;
                    16'h7877: data_out = 8'hEF;
                    16'h7878: data_out = 8'hF0;
                    16'h7879: data_out = 8'hF1;
                    16'h787A: data_out = 8'hF2;
                    16'h787B: data_out = 8'hF3;
                    16'h787C: data_out = 8'hF4;
                    16'h787D: data_out = 8'hF5;
                    16'h787E: data_out = 8'hF6;
                    16'h787F: data_out = 8'hF7;
                    16'h7880: data_out = 8'h78;
                    16'h7881: data_out = 8'h77;
                    16'h7882: data_out = 8'h76;
                    16'h7883: data_out = 8'h75;
                    16'h7884: data_out = 8'h74;
                    16'h7885: data_out = 8'h73;
                    16'h7886: data_out = 8'h72;
                    16'h7887: data_out = 8'h71;
                    16'h7888: data_out = 8'h70;
                    16'h7889: data_out = 8'h6F;
                    16'h788A: data_out = 8'h6E;
                    16'h788B: data_out = 8'h6D;
                    16'h788C: data_out = 8'h6C;
                    16'h788D: data_out = 8'h6B;
                    16'h788E: data_out = 8'h6A;
                    16'h788F: data_out = 8'h69;
                    16'h7890: data_out = 8'h68;
                    16'h7891: data_out = 8'h67;
                    16'h7892: data_out = 8'h66;
                    16'h7893: data_out = 8'h65;
                    16'h7894: data_out = 8'h64;
                    16'h7895: data_out = 8'h63;
                    16'h7896: data_out = 8'h62;
                    16'h7897: data_out = 8'h61;
                    16'h7898: data_out = 8'h60;
                    16'h7899: data_out = 8'h5F;
                    16'h789A: data_out = 8'h5E;
                    16'h789B: data_out = 8'h5D;
                    16'h789C: data_out = 8'h5C;
                    16'h789D: data_out = 8'h5B;
                    16'h789E: data_out = 8'h5A;
                    16'h789F: data_out = 8'h59;
                    16'h78A0: data_out = 8'h58;
                    16'h78A1: data_out = 8'h57;
                    16'h78A2: data_out = 8'h56;
                    16'h78A3: data_out = 8'h55;
                    16'h78A4: data_out = 8'h54;
                    16'h78A5: data_out = 8'h53;
                    16'h78A6: data_out = 8'h52;
                    16'h78A7: data_out = 8'h51;
                    16'h78A8: data_out = 8'h50;
                    16'h78A9: data_out = 8'h4F;
                    16'h78AA: data_out = 8'h4E;
                    16'h78AB: data_out = 8'h4D;
                    16'h78AC: data_out = 8'h4C;
                    16'h78AD: data_out = 8'h4B;
                    16'h78AE: data_out = 8'h4A;
                    16'h78AF: data_out = 8'h49;
                    16'h78B0: data_out = 8'h48;
                    16'h78B1: data_out = 8'h47;
                    16'h78B2: data_out = 8'h46;
                    16'h78B3: data_out = 8'h45;
                    16'h78B4: data_out = 8'h44;
                    16'h78B5: data_out = 8'h43;
                    16'h78B6: data_out = 8'h42;
                    16'h78B7: data_out = 8'h41;
                    16'h78B8: data_out = 8'h40;
                    16'h78B9: data_out = 8'h3F;
                    16'h78BA: data_out = 8'h3E;
                    16'h78BB: data_out = 8'h3D;
                    16'h78BC: data_out = 8'h3C;
                    16'h78BD: data_out = 8'h3B;
                    16'h78BE: data_out = 8'h3A;
                    16'h78BF: data_out = 8'h39;
                    16'h78C0: data_out = 8'h38;
                    16'h78C1: data_out = 8'h37;
                    16'h78C2: data_out = 8'h36;
                    16'h78C3: data_out = 8'h35;
                    16'h78C4: data_out = 8'h34;
                    16'h78C5: data_out = 8'h33;
                    16'h78C6: data_out = 8'h32;
                    16'h78C7: data_out = 8'h31;
                    16'h78C8: data_out = 8'h30;
                    16'h78C9: data_out = 8'h2F;
                    16'h78CA: data_out = 8'h2E;
                    16'h78CB: data_out = 8'h2D;
                    16'h78CC: data_out = 8'h2C;
                    16'h78CD: data_out = 8'h2B;
                    16'h78CE: data_out = 8'h2A;
                    16'h78CF: data_out = 8'h29;
                    16'h78D0: data_out = 8'h28;
                    16'h78D1: data_out = 8'h27;
                    16'h78D2: data_out = 8'h26;
                    16'h78D3: data_out = 8'h25;
                    16'h78D4: data_out = 8'h24;
                    16'h78D5: data_out = 8'h23;
                    16'h78D6: data_out = 8'h22;
                    16'h78D7: data_out = 8'h21;
                    16'h78D8: data_out = 8'h20;
                    16'h78D9: data_out = 8'h1F;
                    16'h78DA: data_out = 8'h1E;
                    16'h78DB: data_out = 8'h1D;
                    16'h78DC: data_out = 8'h1C;
                    16'h78DD: data_out = 8'h1B;
                    16'h78DE: data_out = 8'h1A;
                    16'h78DF: data_out = 8'h19;
                    16'h78E0: data_out = 8'h18;
                    16'h78E1: data_out = 8'h17;
                    16'h78E2: data_out = 8'h16;
                    16'h78E3: data_out = 8'h15;
                    16'h78E4: data_out = 8'h14;
                    16'h78E5: data_out = 8'h13;
                    16'h78E6: data_out = 8'h12;
                    16'h78E7: data_out = 8'h11;
                    16'h78E8: data_out = 8'h10;
                    16'h78E9: data_out = 8'hF;
                    16'h78EA: data_out = 8'hE;
                    16'h78EB: data_out = 8'hD;
                    16'h78EC: data_out = 8'hC;
                    16'h78ED: data_out = 8'hB;
                    16'h78EE: data_out = 8'hA;
                    16'h78EF: data_out = 8'h9;
                    16'h78F0: data_out = 8'h8;
                    16'h78F1: data_out = 8'h7;
                    16'h78F2: data_out = 8'h6;
                    16'h78F3: data_out = 8'h5;
                    16'h78F4: data_out = 8'h4;
                    16'h78F5: data_out = 8'h3;
                    16'h78F6: data_out = 8'h2;
                    16'h78F7: data_out = 8'h1;
                    16'h78F8: data_out = 8'h0;
                    16'h78F9: data_out = 8'h81;
                    16'h78FA: data_out = 8'h82;
                    16'h78FB: data_out = 8'h83;
                    16'h78FC: data_out = 8'h84;
                    16'h78FD: data_out = 8'h85;
                    16'h78FE: data_out = 8'h86;
                    16'h78FF: data_out = 8'h87;
                    16'h7900: data_out = 8'h79;
                    16'h7901: data_out = 8'h7A;
                    16'h7902: data_out = 8'h7B;
                    16'h7903: data_out = 8'h7C;
                    16'h7904: data_out = 8'h7D;
                    16'h7905: data_out = 8'h7E;
                    16'h7906: data_out = 8'h7F;
                    16'h7907: data_out = 8'h80;
                    16'h7908: data_out = 8'h81;
                    16'h7909: data_out = 8'h82;
                    16'h790A: data_out = 8'h83;
                    16'h790B: data_out = 8'h84;
                    16'h790C: data_out = 8'h85;
                    16'h790D: data_out = 8'h86;
                    16'h790E: data_out = 8'h87;
                    16'h790F: data_out = 8'h88;
                    16'h7910: data_out = 8'h89;
                    16'h7911: data_out = 8'h8A;
                    16'h7912: data_out = 8'h8B;
                    16'h7913: data_out = 8'h8C;
                    16'h7914: data_out = 8'h8D;
                    16'h7915: data_out = 8'h8E;
                    16'h7916: data_out = 8'h8F;
                    16'h7917: data_out = 8'h90;
                    16'h7918: data_out = 8'h91;
                    16'h7919: data_out = 8'h92;
                    16'h791A: data_out = 8'h93;
                    16'h791B: data_out = 8'h94;
                    16'h791C: data_out = 8'h95;
                    16'h791D: data_out = 8'h96;
                    16'h791E: data_out = 8'h97;
                    16'h791F: data_out = 8'h98;
                    16'h7920: data_out = 8'h99;
                    16'h7921: data_out = 8'h9A;
                    16'h7922: data_out = 8'h9B;
                    16'h7923: data_out = 8'h9C;
                    16'h7924: data_out = 8'h9D;
                    16'h7925: data_out = 8'h9E;
                    16'h7926: data_out = 8'h9F;
                    16'h7927: data_out = 8'hA0;
                    16'h7928: data_out = 8'hA1;
                    16'h7929: data_out = 8'hA2;
                    16'h792A: data_out = 8'hA3;
                    16'h792B: data_out = 8'hA4;
                    16'h792C: data_out = 8'hA5;
                    16'h792D: data_out = 8'hA6;
                    16'h792E: data_out = 8'hA7;
                    16'h792F: data_out = 8'hA8;
                    16'h7930: data_out = 8'hA9;
                    16'h7931: data_out = 8'hAA;
                    16'h7932: data_out = 8'hAB;
                    16'h7933: data_out = 8'hAC;
                    16'h7934: data_out = 8'hAD;
                    16'h7935: data_out = 8'hAE;
                    16'h7936: data_out = 8'hAF;
                    16'h7937: data_out = 8'hB0;
                    16'h7938: data_out = 8'hB1;
                    16'h7939: data_out = 8'hB2;
                    16'h793A: data_out = 8'hB3;
                    16'h793B: data_out = 8'hB4;
                    16'h793C: data_out = 8'hB5;
                    16'h793D: data_out = 8'hB6;
                    16'h793E: data_out = 8'hB7;
                    16'h793F: data_out = 8'hB8;
                    16'h7940: data_out = 8'hB9;
                    16'h7941: data_out = 8'hBA;
                    16'h7942: data_out = 8'hBB;
                    16'h7943: data_out = 8'hBC;
                    16'h7944: data_out = 8'hBD;
                    16'h7945: data_out = 8'hBE;
                    16'h7946: data_out = 8'hBF;
                    16'h7947: data_out = 8'hC0;
                    16'h7948: data_out = 8'hC1;
                    16'h7949: data_out = 8'hC2;
                    16'h794A: data_out = 8'hC3;
                    16'h794B: data_out = 8'hC4;
                    16'h794C: data_out = 8'hC5;
                    16'h794D: data_out = 8'hC6;
                    16'h794E: data_out = 8'hC7;
                    16'h794F: data_out = 8'hC8;
                    16'h7950: data_out = 8'hC9;
                    16'h7951: data_out = 8'hCA;
                    16'h7952: data_out = 8'hCB;
                    16'h7953: data_out = 8'hCC;
                    16'h7954: data_out = 8'hCD;
                    16'h7955: data_out = 8'hCE;
                    16'h7956: data_out = 8'hCF;
                    16'h7957: data_out = 8'hD0;
                    16'h7958: data_out = 8'hD1;
                    16'h7959: data_out = 8'hD2;
                    16'h795A: data_out = 8'hD3;
                    16'h795B: data_out = 8'hD4;
                    16'h795C: data_out = 8'hD5;
                    16'h795D: data_out = 8'hD6;
                    16'h795E: data_out = 8'hD7;
                    16'h795F: data_out = 8'hD8;
                    16'h7960: data_out = 8'hD9;
                    16'h7961: data_out = 8'hDA;
                    16'h7962: data_out = 8'hDB;
                    16'h7963: data_out = 8'hDC;
                    16'h7964: data_out = 8'hDD;
                    16'h7965: data_out = 8'hDE;
                    16'h7966: data_out = 8'hDF;
                    16'h7967: data_out = 8'hE0;
                    16'h7968: data_out = 8'hE1;
                    16'h7969: data_out = 8'hE2;
                    16'h796A: data_out = 8'hE3;
                    16'h796B: data_out = 8'hE4;
                    16'h796C: data_out = 8'hE5;
                    16'h796D: data_out = 8'hE6;
                    16'h796E: data_out = 8'hE7;
                    16'h796F: data_out = 8'hE8;
                    16'h7970: data_out = 8'hE9;
                    16'h7971: data_out = 8'hEA;
                    16'h7972: data_out = 8'hEB;
                    16'h7973: data_out = 8'hEC;
                    16'h7974: data_out = 8'hED;
                    16'h7975: data_out = 8'hEE;
                    16'h7976: data_out = 8'hEF;
                    16'h7977: data_out = 8'hF0;
                    16'h7978: data_out = 8'hF1;
                    16'h7979: data_out = 8'hF2;
                    16'h797A: data_out = 8'hF3;
                    16'h797B: data_out = 8'hF4;
                    16'h797C: data_out = 8'hF5;
                    16'h797D: data_out = 8'hF6;
                    16'h797E: data_out = 8'hF7;
                    16'h797F: data_out = 8'hF8;
                    16'h7980: data_out = 8'h79;
                    16'h7981: data_out = 8'h78;
                    16'h7982: data_out = 8'h77;
                    16'h7983: data_out = 8'h76;
                    16'h7984: data_out = 8'h75;
                    16'h7985: data_out = 8'h74;
                    16'h7986: data_out = 8'h73;
                    16'h7987: data_out = 8'h72;
                    16'h7988: data_out = 8'h71;
                    16'h7989: data_out = 8'h70;
                    16'h798A: data_out = 8'h6F;
                    16'h798B: data_out = 8'h6E;
                    16'h798C: data_out = 8'h6D;
                    16'h798D: data_out = 8'h6C;
                    16'h798E: data_out = 8'h6B;
                    16'h798F: data_out = 8'h6A;
                    16'h7990: data_out = 8'h69;
                    16'h7991: data_out = 8'h68;
                    16'h7992: data_out = 8'h67;
                    16'h7993: data_out = 8'h66;
                    16'h7994: data_out = 8'h65;
                    16'h7995: data_out = 8'h64;
                    16'h7996: data_out = 8'h63;
                    16'h7997: data_out = 8'h62;
                    16'h7998: data_out = 8'h61;
                    16'h7999: data_out = 8'h60;
                    16'h799A: data_out = 8'h5F;
                    16'h799B: data_out = 8'h5E;
                    16'h799C: data_out = 8'h5D;
                    16'h799D: data_out = 8'h5C;
                    16'h799E: data_out = 8'h5B;
                    16'h799F: data_out = 8'h5A;
                    16'h79A0: data_out = 8'h59;
                    16'h79A1: data_out = 8'h58;
                    16'h79A2: data_out = 8'h57;
                    16'h79A3: data_out = 8'h56;
                    16'h79A4: data_out = 8'h55;
                    16'h79A5: data_out = 8'h54;
                    16'h79A6: data_out = 8'h53;
                    16'h79A7: data_out = 8'h52;
                    16'h79A8: data_out = 8'h51;
                    16'h79A9: data_out = 8'h50;
                    16'h79AA: data_out = 8'h4F;
                    16'h79AB: data_out = 8'h4E;
                    16'h79AC: data_out = 8'h4D;
                    16'h79AD: data_out = 8'h4C;
                    16'h79AE: data_out = 8'h4B;
                    16'h79AF: data_out = 8'h4A;
                    16'h79B0: data_out = 8'h49;
                    16'h79B1: data_out = 8'h48;
                    16'h79B2: data_out = 8'h47;
                    16'h79B3: data_out = 8'h46;
                    16'h79B4: data_out = 8'h45;
                    16'h79B5: data_out = 8'h44;
                    16'h79B6: data_out = 8'h43;
                    16'h79B7: data_out = 8'h42;
                    16'h79B8: data_out = 8'h41;
                    16'h79B9: data_out = 8'h40;
                    16'h79BA: data_out = 8'h3F;
                    16'h79BB: data_out = 8'h3E;
                    16'h79BC: data_out = 8'h3D;
                    16'h79BD: data_out = 8'h3C;
                    16'h79BE: data_out = 8'h3B;
                    16'h79BF: data_out = 8'h3A;
                    16'h79C0: data_out = 8'h39;
                    16'h79C1: data_out = 8'h38;
                    16'h79C2: data_out = 8'h37;
                    16'h79C3: data_out = 8'h36;
                    16'h79C4: data_out = 8'h35;
                    16'h79C5: data_out = 8'h34;
                    16'h79C6: data_out = 8'h33;
                    16'h79C7: data_out = 8'h32;
                    16'h79C8: data_out = 8'h31;
                    16'h79C9: data_out = 8'h30;
                    16'h79CA: data_out = 8'h2F;
                    16'h79CB: data_out = 8'h2E;
                    16'h79CC: data_out = 8'h2D;
                    16'h79CD: data_out = 8'h2C;
                    16'h79CE: data_out = 8'h2B;
                    16'h79CF: data_out = 8'h2A;
                    16'h79D0: data_out = 8'h29;
                    16'h79D1: data_out = 8'h28;
                    16'h79D2: data_out = 8'h27;
                    16'h79D3: data_out = 8'h26;
                    16'h79D4: data_out = 8'h25;
                    16'h79D5: data_out = 8'h24;
                    16'h79D6: data_out = 8'h23;
                    16'h79D7: data_out = 8'h22;
                    16'h79D8: data_out = 8'h21;
                    16'h79D9: data_out = 8'h20;
                    16'h79DA: data_out = 8'h1F;
                    16'h79DB: data_out = 8'h1E;
                    16'h79DC: data_out = 8'h1D;
                    16'h79DD: data_out = 8'h1C;
                    16'h79DE: data_out = 8'h1B;
                    16'h79DF: data_out = 8'h1A;
                    16'h79E0: data_out = 8'h19;
                    16'h79E1: data_out = 8'h18;
                    16'h79E2: data_out = 8'h17;
                    16'h79E3: data_out = 8'h16;
                    16'h79E4: data_out = 8'h15;
                    16'h79E5: data_out = 8'h14;
                    16'h79E6: data_out = 8'h13;
                    16'h79E7: data_out = 8'h12;
                    16'h79E8: data_out = 8'h11;
                    16'h79E9: data_out = 8'h10;
                    16'h79EA: data_out = 8'hF;
                    16'h79EB: data_out = 8'hE;
                    16'h79EC: data_out = 8'hD;
                    16'h79ED: data_out = 8'hC;
                    16'h79EE: data_out = 8'hB;
                    16'h79EF: data_out = 8'hA;
                    16'h79F0: data_out = 8'h9;
                    16'h79F1: data_out = 8'h8;
                    16'h79F2: data_out = 8'h7;
                    16'h79F3: data_out = 8'h6;
                    16'h79F4: data_out = 8'h5;
                    16'h79F5: data_out = 8'h4;
                    16'h79F6: data_out = 8'h3;
                    16'h79F7: data_out = 8'h2;
                    16'h79F8: data_out = 8'h1;
                    16'h79F9: data_out = 8'h0;
                    16'h79FA: data_out = 8'h81;
                    16'h79FB: data_out = 8'h82;
                    16'h79FC: data_out = 8'h83;
                    16'h79FD: data_out = 8'h84;
                    16'h79FE: data_out = 8'h85;
                    16'h79FF: data_out = 8'h86;
                    16'h7A00: data_out = 8'h7A;
                    16'h7A01: data_out = 8'h7B;
                    16'h7A02: data_out = 8'h7C;
                    16'h7A03: data_out = 8'h7D;
                    16'h7A04: data_out = 8'h7E;
                    16'h7A05: data_out = 8'h7F;
                    16'h7A06: data_out = 8'h80;
                    16'h7A07: data_out = 8'h81;
                    16'h7A08: data_out = 8'h82;
                    16'h7A09: data_out = 8'h83;
                    16'h7A0A: data_out = 8'h84;
                    16'h7A0B: data_out = 8'h85;
                    16'h7A0C: data_out = 8'h86;
                    16'h7A0D: data_out = 8'h87;
                    16'h7A0E: data_out = 8'h88;
                    16'h7A0F: data_out = 8'h89;
                    16'h7A10: data_out = 8'h8A;
                    16'h7A11: data_out = 8'h8B;
                    16'h7A12: data_out = 8'h8C;
                    16'h7A13: data_out = 8'h8D;
                    16'h7A14: data_out = 8'h8E;
                    16'h7A15: data_out = 8'h8F;
                    16'h7A16: data_out = 8'h90;
                    16'h7A17: data_out = 8'h91;
                    16'h7A18: data_out = 8'h92;
                    16'h7A19: data_out = 8'h93;
                    16'h7A1A: data_out = 8'h94;
                    16'h7A1B: data_out = 8'h95;
                    16'h7A1C: data_out = 8'h96;
                    16'h7A1D: data_out = 8'h97;
                    16'h7A1E: data_out = 8'h98;
                    16'h7A1F: data_out = 8'h99;
                    16'h7A20: data_out = 8'h9A;
                    16'h7A21: data_out = 8'h9B;
                    16'h7A22: data_out = 8'h9C;
                    16'h7A23: data_out = 8'h9D;
                    16'h7A24: data_out = 8'h9E;
                    16'h7A25: data_out = 8'h9F;
                    16'h7A26: data_out = 8'hA0;
                    16'h7A27: data_out = 8'hA1;
                    16'h7A28: data_out = 8'hA2;
                    16'h7A29: data_out = 8'hA3;
                    16'h7A2A: data_out = 8'hA4;
                    16'h7A2B: data_out = 8'hA5;
                    16'h7A2C: data_out = 8'hA6;
                    16'h7A2D: data_out = 8'hA7;
                    16'h7A2E: data_out = 8'hA8;
                    16'h7A2F: data_out = 8'hA9;
                    16'h7A30: data_out = 8'hAA;
                    16'h7A31: data_out = 8'hAB;
                    16'h7A32: data_out = 8'hAC;
                    16'h7A33: data_out = 8'hAD;
                    16'h7A34: data_out = 8'hAE;
                    16'h7A35: data_out = 8'hAF;
                    16'h7A36: data_out = 8'hB0;
                    16'h7A37: data_out = 8'hB1;
                    16'h7A38: data_out = 8'hB2;
                    16'h7A39: data_out = 8'hB3;
                    16'h7A3A: data_out = 8'hB4;
                    16'h7A3B: data_out = 8'hB5;
                    16'h7A3C: data_out = 8'hB6;
                    16'h7A3D: data_out = 8'hB7;
                    16'h7A3E: data_out = 8'hB8;
                    16'h7A3F: data_out = 8'hB9;
                    16'h7A40: data_out = 8'hBA;
                    16'h7A41: data_out = 8'hBB;
                    16'h7A42: data_out = 8'hBC;
                    16'h7A43: data_out = 8'hBD;
                    16'h7A44: data_out = 8'hBE;
                    16'h7A45: data_out = 8'hBF;
                    16'h7A46: data_out = 8'hC0;
                    16'h7A47: data_out = 8'hC1;
                    16'h7A48: data_out = 8'hC2;
                    16'h7A49: data_out = 8'hC3;
                    16'h7A4A: data_out = 8'hC4;
                    16'h7A4B: data_out = 8'hC5;
                    16'h7A4C: data_out = 8'hC6;
                    16'h7A4D: data_out = 8'hC7;
                    16'h7A4E: data_out = 8'hC8;
                    16'h7A4F: data_out = 8'hC9;
                    16'h7A50: data_out = 8'hCA;
                    16'h7A51: data_out = 8'hCB;
                    16'h7A52: data_out = 8'hCC;
                    16'h7A53: data_out = 8'hCD;
                    16'h7A54: data_out = 8'hCE;
                    16'h7A55: data_out = 8'hCF;
                    16'h7A56: data_out = 8'hD0;
                    16'h7A57: data_out = 8'hD1;
                    16'h7A58: data_out = 8'hD2;
                    16'h7A59: data_out = 8'hD3;
                    16'h7A5A: data_out = 8'hD4;
                    16'h7A5B: data_out = 8'hD5;
                    16'h7A5C: data_out = 8'hD6;
                    16'h7A5D: data_out = 8'hD7;
                    16'h7A5E: data_out = 8'hD8;
                    16'h7A5F: data_out = 8'hD9;
                    16'h7A60: data_out = 8'hDA;
                    16'h7A61: data_out = 8'hDB;
                    16'h7A62: data_out = 8'hDC;
                    16'h7A63: data_out = 8'hDD;
                    16'h7A64: data_out = 8'hDE;
                    16'h7A65: data_out = 8'hDF;
                    16'h7A66: data_out = 8'hE0;
                    16'h7A67: data_out = 8'hE1;
                    16'h7A68: data_out = 8'hE2;
                    16'h7A69: data_out = 8'hE3;
                    16'h7A6A: data_out = 8'hE4;
                    16'h7A6B: data_out = 8'hE5;
                    16'h7A6C: data_out = 8'hE6;
                    16'h7A6D: data_out = 8'hE7;
                    16'h7A6E: data_out = 8'hE8;
                    16'h7A6F: data_out = 8'hE9;
                    16'h7A70: data_out = 8'hEA;
                    16'h7A71: data_out = 8'hEB;
                    16'h7A72: data_out = 8'hEC;
                    16'h7A73: data_out = 8'hED;
                    16'h7A74: data_out = 8'hEE;
                    16'h7A75: data_out = 8'hEF;
                    16'h7A76: data_out = 8'hF0;
                    16'h7A77: data_out = 8'hF1;
                    16'h7A78: data_out = 8'hF2;
                    16'h7A79: data_out = 8'hF3;
                    16'h7A7A: data_out = 8'hF4;
                    16'h7A7B: data_out = 8'hF5;
                    16'h7A7C: data_out = 8'hF6;
                    16'h7A7D: data_out = 8'hF7;
                    16'h7A7E: data_out = 8'hF8;
                    16'h7A7F: data_out = 8'hF9;
                    16'h7A80: data_out = 8'h7A;
                    16'h7A81: data_out = 8'h79;
                    16'h7A82: data_out = 8'h78;
                    16'h7A83: data_out = 8'h77;
                    16'h7A84: data_out = 8'h76;
                    16'h7A85: data_out = 8'h75;
                    16'h7A86: data_out = 8'h74;
                    16'h7A87: data_out = 8'h73;
                    16'h7A88: data_out = 8'h72;
                    16'h7A89: data_out = 8'h71;
                    16'h7A8A: data_out = 8'h70;
                    16'h7A8B: data_out = 8'h6F;
                    16'h7A8C: data_out = 8'h6E;
                    16'h7A8D: data_out = 8'h6D;
                    16'h7A8E: data_out = 8'h6C;
                    16'h7A8F: data_out = 8'h6B;
                    16'h7A90: data_out = 8'h6A;
                    16'h7A91: data_out = 8'h69;
                    16'h7A92: data_out = 8'h68;
                    16'h7A93: data_out = 8'h67;
                    16'h7A94: data_out = 8'h66;
                    16'h7A95: data_out = 8'h65;
                    16'h7A96: data_out = 8'h64;
                    16'h7A97: data_out = 8'h63;
                    16'h7A98: data_out = 8'h62;
                    16'h7A99: data_out = 8'h61;
                    16'h7A9A: data_out = 8'h60;
                    16'h7A9B: data_out = 8'h5F;
                    16'h7A9C: data_out = 8'h5E;
                    16'h7A9D: data_out = 8'h5D;
                    16'h7A9E: data_out = 8'h5C;
                    16'h7A9F: data_out = 8'h5B;
                    16'h7AA0: data_out = 8'h5A;
                    16'h7AA1: data_out = 8'h59;
                    16'h7AA2: data_out = 8'h58;
                    16'h7AA3: data_out = 8'h57;
                    16'h7AA4: data_out = 8'h56;
                    16'h7AA5: data_out = 8'h55;
                    16'h7AA6: data_out = 8'h54;
                    16'h7AA7: data_out = 8'h53;
                    16'h7AA8: data_out = 8'h52;
                    16'h7AA9: data_out = 8'h51;
                    16'h7AAA: data_out = 8'h50;
                    16'h7AAB: data_out = 8'h4F;
                    16'h7AAC: data_out = 8'h4E;
                    16'h7AAD: data_out = 8'h4D;
                    16'h7AAE: data_out = 8'h4C;
                    16'h7AAF: data_out = 8'h4B;
                    16'h7AB0: data_out = 8'h4A;
                    16'h7AB1: data_out = 8'h49;
                    16'h7AB2: data_out = 8'h48;
                    16'h7AB3: data_out = 8'h47;
                    16'h7AB4: data_out = 8'h46;
                    16'h7AB5: data_out = 8'h45;
                    16'h7AB6: data_out = 8'h44;
                    16'h7AB7: data_out = 8'h43;
                    16'h7AB8: data_out = 8'h42;
                    16'h7AB9: data_out = 8'h41;
                    16'h7ABA: data_out = 8'h40;
                    16'h7ABB: data_out = 8'h3F;
                    16'h7ABC: data_out = 8'h3E;
                    16'h7ABD: data_out = 8'h3D;
                    16'h7ABE: data_out = 8'h3C;
                    16'h7ABF: data_out = 8'h3B;
                    16'h7AC0: data_out = 8'h3A;
                    16'h7AC1: data_out = 8'h39;
                    16'h7AC2: data_out = 8'h38;
                    16'h7AC3: data_out = 8'h37;
                    16'h7AC4: data_out = 8'h36;
                    16'h7AC5: data_out = 8'h35;
                    16'h7AC6: data_out = 8'h34;
                    16'h7AC7: data_out = 8'h33;
                    16'h7AC8: data_out = 8'h32;
                    16'h7AC9: data_out = 8'h31;
                    16'h7ACA: data_out = 8'h30;
                    16'h7ACB: data_out = 8'h2F;
                    16'h7ACC: data_out = 8'h2E;
                    16'h7ACD: data_out = 8'h2D;
                    16'h7ACE: data_out = 8'h2C;
                    16'h7ACF: data_out = 8'h2B;
                    16'h7AD0: data_out = 8'h2A;
                    16'h7AD1: data_out = 8'h29;
                    16'h7AD2: data_out = 8'h28;
                    16'h7AD3: data_out = 8'h27;
                    16'h7AD4: data_out = 8'h26;
                    16'h7AD5: data_out = 8'h25;
                    16'h7AD6: data_out = 8'h24;
                    16'h7AD7: data_out = 8'h23;
                    16'h7AD8: data_out = 8'h22;
                    16'h7AD9: data_out = 8'h21;
                    16'h7ADA: data_out = 8'h20;
                    16'h7ADB: data_out = 8'h1F;
                    16'h7ADC: data_out = 8'h1E;
                    16'h7ADD: data_out = 8'h1D;
                    16'h7ADE: data_out = 8'h1C;
                    16'h7ADF: data_out = 8'h1B;
                    16'h7AE0: data_out = 8'h1A;
                    16'h7AE1: data_out = 8'h19;
                    16'h7AE2: data_out = 8'h18;
                    16'h7AE3: data_out = 8'h17;
                    16'h7AE4: data_out = 8'h16;
                    16'h7AE5: data_out = 8'h15;
                    16'h7AE6: data_out = 8'h14;
                    16'h7AE7: data_out = 8'h13;
                    16'h7AE8: data_out = 8'h12;
                    16'h7AE9: data_out = 8'h11;
                    16'h7AEA: data_out = 8'h10;
                    16'h7AEB: data_out = 8'hF;
                    16'h7AEC: data_out = 8'hE;
                    16'h7AED: data_out = 8'hD;
                    16'h7AEE: data_out = 8'hC;
                    16'h7AEF: data_out = 8'hB;
                    16'h7AF0: data_out = 8'hA;
                    16'h7AF1: data_out = 8'h9;
                    16'h7AF2: data_out = 8'h8;
                    16'h7AF3: data_out = 8'h7;
                    16'h7AF4: data_out = 8'h6;
                    16'h7AF5: data_out = 8'h5;
                    16'h7AF6: data_out = 8'h4;
                    16'h7AF7: data_out = 8'h3;
                    16'h7AF8: data_out = 8'h2;
                    16'h7AF9: data_out = 8'h1;
                    16'h7AFA: data_out = 8'h0;
                    16'h7AFB: data_out = 8'h81;
                    16'h7AFC: data_out = 8'h82;
                    16'h7AFD: data_out = 8'h83;
                    16'h7AFE: data_out = 8'h84;
                    16'h7AFF: data_out = 8'h85;
                    16'h7B00: data_out = 8'h7B;
                    16'h7B01: data_out = 8'h7C;
                    16'h7B02: data_out = 8'h7D;
                    16'h7B03: data_out = 8'h7E;
                    16'h7B04: data_out = 8'h7F;
                    16'h7B05: data_out = 8'h80;
                    16'h7B06: data_out = 8'h81;
                    16'h7B07: data_out = 8'h82;
                    16'h7B08: data_out = 8'h83;
                    16'h7B09: data_out = 8'h84;
                    16'h7B0A: data_out = 8'h85;
                    16'h7B0B: data_out = 8'h86;
                    16'h7B0C: data_out = 8'h87;
                    16'h7B0D: data_out = 8'h88;
                    16'h7B0E: data_out = 8'h89;
                    16'h7B0F: data_out = 8'h8A;
                    16'h7B10: data_out = 8'h8B;
                    16'h7B11: data_out = 8'h8C;
                    16'h7B12: data_out = 8'h8D;
                    16'h7B13: data_out = 8'h8E;
                    16'h7B14: data_out = 8'h8F;
                    16'h7B15: data_out = 8'h90;
                    16'h7B16: data_out = 8'h91;
                    16'h7B17: data_out = 8'h92;
                    16'h7B18: data_out = 8'h93;
                    16'h7B19: data_out = 8'h94;
                    16'h7B1A: data_out = 8'h95;
                    16'h7B1B: data_out = 8'h96;
                    16'h7B1C: data_out = 8'h97;
                    16'h7B1D: data_out = 8'h98;
                    16'h7B1E: data_out = 8'h99;
                    16'h7B1F: data_out = 8'h9A;
                    16'h7B20: data_out = 8'h9B;
                    16'h7B21: data_out = 8'h9C;
                    16'h7B22: data_out = 8'h9D;
                    16'h7B23: data_out = 8'h9E;
                    16'h7B24: data_out = 8'h9F;
                    16'h7B25: data_out = 8'hA0;
                    16'h7B26: data_out = 8'hA1;
                    16'h7B27: data_out = 8'hA2;
                    16'h7B28: data_out = 8'hA3;
                    16'h7B29: data_out = 8'hA4;
                    16'h7B2A: data_out = 8'hA5;
                    16'h7B2B: data_out = 8'hA6;
                    16'h7B2C: data_out = 8'hA7;
                    16'h7B2D: data_out = 8'hA8;
                    16'h7B2E: data_out = 8'hA9;
                    16'h7B2F: data_out = 8'hAA;
                    16'h7B30: data_out = 8'hAB;
                    16'h7B31: data_out = 8'hAC;
                    16'h7B32: data_out = 8'hAD;
                    16'h7B33: data_out = 8'hAE;
                    16'h7B34: data_out = 8'hAF;
                    16'h7B35: data_out = 8'hB0;
                    16'h7B36: data_out = 8'hB1;
                    16'h7B37: data_out = 8'hB2;
                    16'h7B38: data_out = 8'hB3;
                    16'h7B39: data_out = 8'hB4;
                    16'h7B3A: data_out = 8'hB5;
                    16'h7B3B: data_out = 8'hB6;
                    16'h7B3C: data_out = 8'hB7;
                    16'h7B3D: data_out = 8'hB8;
                    16'h7B3E: data_out = 8'hB9;
                    16'h7B3F: data_out = 8'hBA;
                    16'h7B40: data_out = 8'hBB;
                    16'h7B41: data_out = 8'hBC;
                    16'h7B42: data_out = 8'hBD;
                    16'h7B43: data_out = 8'hBE;
                    16'h7B44: data_out = 8'hBF;
                    16'h7B45: data_out = 8'hC0;
                    16'h7B46: data_out = 8'hC1;
                    16'h7B47: data_out = 8'hC2;
                    16'h7B48: data_out = 8'hC3;
                    16'h7B49: data_out = 8'hC4;
                    16'h7B4A: data_out = 8'hC5;
                    16'h7B4B: data_out = 8'hC6;
                    16'h7B4C: data_out = 8'hC7;
                    16'h7B4D: data_out = 8'hC8;
                    16'h7B4E: data_out = 8'hC9;
                    16'h7B4F: data_out = 8'hCA;
                    16'h7B50: data_out = 8'hCB;
                    16'h7B51: data_out = 8'hCC;
                    16'h7B52: data_out = 8'hCD;
                    16'h7B53: data_out = 8'hCE;
                    16'h7B54: data_out = 8'hCF;
                    16'h7B55: data_out = 8'hD0;
                    16'h7B56: data_out = 8'hD1;
                    16'h7B57: data_out = 8'hD2;
                    16'h7B58: data_out = 8'hD3;
                    16'h7B59: data_out = 8'hD4;
                    16'h7B5A: data_out = 8'hD5;
                    16'h7B5B: data_out = 8'hD6;
                    16'h7B5C: data_out = 8'hD7;
                    16'h7B5D: data_out = 8'hD8;
                    16'h7B5E: data_out = 8'hD9;
                    16'h7B5F: data_out = 8'hDA;
                    16'h7B60: data_out = 8'hDB;
                    16'h7B61: data_out = 8'hDC;
                    16'h7B62: data_out = 8'hDD;
                    16'h7B63: data_out = 8'hDE;
                    16'h7B64: data_out = 8'hDF;
                    16'h7B65: data_out = 8'hE0;
                    16'h7B66: data_out = 8'hE1;
                    16'h7B67: data_out = 8'hE2;
                    16'h7B68: data_out = 8'hE3;
                    16'h7B69: data_out = 8'hE4;
                    16'h7B6A: data_out = 8'hE5;
                    16'h7B6B: data_out = 8'hE6;
                    16'h7B6C: data_out = 8'hE7;
                    16'h7B6D: data_out = 8'hE8;
                    16'h7B6E: data_out = 8'hE9;
                    16'h7B6F: data_out = 8'hEA;
                    16'h7B70: data_out = 8'hEB;
                    16'h7B71: data_out = 8'hEC;
                    16'h7B72: data_out = 8'hED;
                    16'h7B73: data_out = 8'hEE;
                    16'h7B74: data_out = 8'hEF;
                    16'h7B75: data_out = 8'hF0;
                    16'h7B76: data_out = 8'hF1;
                    16'h7B77: data_out = 8'hF2;
                    16'h7B78: data_out = 8'hF3;
                    16'h7B79: data_out = 8'hF4;
                    16'h7B7A: data_out = 8'hF5;
                    16'h7B7B: data_out = 8'hF6;
                    16'h7B7C: data_out = 8'hF7;
                    16'h7B7D: data_out = 8'hF8;
                    16'h7B7E: data_out = 8'hF9;
                    16'h7B7F: data_out = 8'hFA;
                    16'h7B80: data_out = 8'h7B;
                    16'h7B81: data_out = 8'h7A;
                    16'h7B82: data_out = 8'h79;
                    16'h7B83: data_out = 8'h78;
                    16'h7B84: data_out = 8'h77;
                    16'h7B85: data_out = 8'h76;
                    16'h7B86: data_out = 8'h75;
                    16'h7B87: data_out = 8'h74;
                    16'h7B88: data_out = 8'h73;
                    16'h7B89: data_out = 8'h72;
                    16'h7B8A: data_out = 8'h71;
                    16'h7B8B: data_out = 8'h70;
                    16'h7B8C: data_out = 8'h6F;
                    16'h7B8D: data_out = 8'h6E;
                    16'h7B8E: data_out = 8'h6D;
                    16'h7B8F: data_out = 8'h6C;
                    16'h7B90: data_out = 8'h6B;
                    16'h7B91: data_out = 8'h6A;
                    16'h7B92: data_out = 8'h69;
                    16'h7B93: data_out = 8'h68;
                    16'h7B94: data_out = 8'h67;
                    16'h7B95: data_out = 8'h66;
                    16'h7B96: data_out = 8'h65;
                    16'h7B97: data_out = 8'h64;
                    16'h7B98: data_out = 8'h63;
                    16'h7B99: data_out = 8'h62;
                    16'h7B9A: data_out = 8'h61;
                    16'h7B9B: data_out = 8'h60;
                    16'h7B9C: data_out = 8'h5F;
                    16'h7B9D: data_out = 8'h5E;
                    16'h7B9E: data_out = 8'h5D;
                    16'h7B9F: data_out = 8'h5C;
                    16'h7BA0: data_out = 8'h5B;
                    16'h7BA1: data_out = 8'h5A;
                    16'h7BA2: data_out = 8'h59;
                    16'h7BA3: data_out = 8'h58;
                    16'h7BA4: data_out = 8'h57;
                    16'h7BA5: data_out = 8'h56;
                    16'h7BA6: data_out = 8'h55;
                    16'h7BA7: data_out = 8'h54;
                    16'h7BA8: data_out = 8'h53;
                    16'h7BA9: data_out = 8'h52;
                    16'h7BAA: data_out = 8'h51;
                    16'h7BAB: data_out = 8'h50;
                    16'h7BAC: data_out = 8'h4F;
                    16'h7BAD: data_out = 8'h4E;
                    16'h7BAE: data_out = 8'h4D;
                    16'h7BAF: data_out = 8'h4C;
                    16'h7BB0: data_out = 8'h4B;
                    16'h7BB1: data_out = 8'h4A;
                    16'h7BB2: data_out = 8'h49;
                    16'h7BB3: data_out = 8'h48;
                    16'h7BB4: data_out = 8'h47;
                    16'h7BB5: data_out = 8'h46;
                    16'h7BB6: data_out = 8'h45;
                    16'h7BB7: data_out = 8'h44;
                    16'h7BB8: data_out = 8'h43;
                    16'h7BB9: data_out = 8'h42;
                    16'h7BBA: data_out = 8'h41;
                    16'h7BBB: data_out = 8'h40;
                    16'h7BBC: data_out = 8'h3F;
                    16'h7BBD: data_out = 8'h3E;
                    16'h7BBE: data_out = 8'h3D;
                    16'h7BBF: data_out = 8'h3C;
                    16'h7BC0: data_out = 8'h3B;
                    16'h7BC1: data_out = 8'h3A;
                    16'h7BC2: data_out = 8'h39;
                    16'h7BC3: data_out = 8'h38;
                    16'h7BC4: data_out = 8'h37;
                    16'h7BC5: data_out = 8'h36;
                    16'h7BC6: data_out = 8'h35;
                    16'h7BC7: data_out = 8'h34;
                    16'h7BC8: data_out = 8'h33;
                    16'h7BC9: data_out = 8'h32;
                    16'h7BCA: data_out = 8'h31;
                    16'h7BCB: data_out = 8'h30;
                    16'h7BCC: data_out = 8'h2F;
                    16'h7BCD: data_out = 8'h2E;
                    16'h7BCE: data_out = 8'h2D;
                    16'h7BCF: data_out = 8'h2C;
                    16'h7BD0: data_out = 8'h2B;
                    16'h7BD1: data_out = 8'h2A;
                    16'h7BD2: data_out = 8'h29;
                    16'h7BD3: data_out = 8'h28;
                    16'h7BD4: data_out = 8'h27;
                    16'h7BD5: data_out = 8'h26;
                    16'h7BD6: data_out = 8'h25;
                    16'h7BD7: data_out = 8'h24;
                    16'h7BD8: data_out = 8'h23;
                    16'h7BD9: data_out = 8'h22;
                    16'h7BDA: data_out = 8'h21;
                    16'h7BDB: data_out = 8'h20;
                    16'h7BDC: data_out = 8'h1F;
                    16'h7BDD: data_out = 8'h1E;
                    16'h7BDE: data_out = 8'h1D;
                    16'h7BDF: data_out = 8'h1C;
                    16'h7BE0: data_out = 8'h1B;
                    16'h7BE1: data_out = 8'h1A;
                    16'h7BE2: data_out = 8'h19;
                    16'h7BE3: data_out = 8'h18;
                    16'h7BE4: data_out = 8'h17;
                    16'h7BE5: data_out = 8'h16;
                    16'h7BE6: data_out = 8'h15;
                    16'h7BE7: data_out = 8'h14;
                    16'h7BE8: data_out = 8'h13;
                    16'h7BE9: data_out = 8'h12;
                    16'h7BEA: data_out = 8'h11;
                    16'h7BEB: data_out = 8'h10;
                    16'h7BEC: data_out = 8'hF;
                    16'h7BED: data_out = 8'hE;
                    16'h7BEE: data_out = 8'hD;
                    16'h7BEF: data_out = 8'hC;
                    16'h7BF0: data_out = 8'hB;
                    16'h7BF1: data_out = 8'hA;
                    16'h7BF2: data_out = 8'h9;
                    16'h7BF3: data_out = 8'h8;
                    16'h7BF4: data_out = 8'h7;
                    16'h7BF5: data_out = 8'h6;
                    16'h7BF6: data_out = 8'h5;
                    16'h7BF7: data_out = 8'h4;
                    16'h7BF8: data_out = 8'h3;
                    16'h7BF9: data_out = 8'h2;
                    16'h7BFA: data_out = 8'h1;
                    16'h7BFB: data_out = 8'h0;
                    16'h7BFC: data_out = 8'h81;
                    16'h7BFD: data_out = 8'h82;
                    16'h7BFE: data_out = 8'h83;
                    16'h7BFF: data_out = 8'h84;
                    16'h7C00: data_out = 8'h7C;
                    16'h7C01: data_out = 8'h7D;
                    16'h7C02: data_out = 8'h7E;
                    16'h7C03: data_out = 8'h7F;
                    16'h7C04: data_out = 8'h80;
                    16'h7C05: data_out = 8'h81;
                    16'h7C06: data_out = 8'h82;
                    16'h7C07: data_out = 8'h83;
                    16'h7C08: data_out = 8'h84;
                    16'h7C09: data_out = 8'h85;
                    16'h7C0A: data_out = 8'h86;
                    16'h7C0B: data_out = 8'h87;
                    16'h7C0C: data_out = 8'h88;
                    16'h7C0D: data_out = 8'h89;
                    16'h7C0E: data_out = 8'h8A;
                    16'h7C0F: data_out = 8'h8B;
                    16'h7C10: data_out = 8'h8C;
                    16'h7C11: data_out = 8'h8D;
                    16'h7C12: data_out = 8'h8E;
                    16'h7C13: data_out = 8'h8F;
                    16'h7C14: data_out = 8'h90;
                    16'h7C15: data_out = 8'h91;
                    16'h7C16: data_out = 8'h92;
                    16'h7C17: data_out = 8'h93;
                    16'h7C18: data_out = 8'h94;
                    16'h7C19: data_out = 8'h95;
                    16'h7C1A: data_out = 8'h96;
                    16'h7C1B: data_out = 8'h97;
                    16'h7C1C: data_out = 8'h98;
                    16'h7C1D: data_out = 8'h99;
                    16'h7C1E: data_out = 8'h9A;
                    16'h7C1F: data_out = 8'h9B;
                    16'h7C20: data_out = 8'h9C;
                    16'h7C21: data_out = 8'h9D;
                    16'h7C22: data_out = 8'h9E;
                    16'h7C23: data_out = 8'h9F;
                    16'h7C24: data_out = 8'hA0;
                    16'h7C25: data_out = 8'hA1;
                    16'h7C26: data_out = 8'hA2;
                    16'h7C27: data_out = 8'hA3;
                    16'h7C28: data_out = 8'hA4;
                    16'h7C29: data_out = 8'hA5;
                    16'h7C2A: data_out = 8'hA6;
                    16'h7C2B: data_out = 8'hA7;
                    16'h7C2C: data_out = 8'hA8;
                    16'h7C2D: data_out = 8'hA9;
                    16'h7C2E: data_out = 8'hAA;
                    16'h7C2F: data_out = 8'hAB;
                    16'h7C30: data_out = 8'hAC;
                    16'h7C31: data_out = 8'hAD;
                    16'h7C32: data_out = 8'hAE;
                    16'h7C33: data_out = 8'hAF;
                    16'h7C34: data_out = 8'hB0;
                    16'h7C35: data_out = 8'hB1;
                    16'h7C36: data_out = 8'hB2;
                    16'h7C37: data_out = 8'hB3;
                    16'h7C38: data_out = 8'hB4;
                    16'h7C39: data_out = 8'hB5;
                    16'h7C3A: data_out = 8'hB6;
                    16'h7C3B: data_out = 8'hB7;
                    16'h7C3C: data_out = 8'hB8;
                    16'h7C3D: data_out = 8'hB9;
                    16'h7C3E: data_out = 8'hBA;
                    16'h7C3F: data_out = 8'hBB;
                    16'h7C40: data_out = 8'hBC;
                    16'h7C41: data_out = 8'hBD;
                    16'h7C42: data_out = 8'hBE;
                    16'h7C43: data_out = 8'hBF;
                    16'h7C44: data_out = 8'hC0;
                    16'h7C45: data_out = 8'hC1;
                    16'h7C46: data_out = 8'hC2;
                    16'h7C47: data_out = 8'hC3;
                    16'h7C48: data_out = 8'hC4;
                    16'h7C49: data_out = 8'hC5;
                    16'h7C4A: data_out = 8'hC6;
                    16'h7C4B: data_out = 8'hC7;
                    16'h7C4C: data_out = 8'hC8;
                    16'h7C4D: data_out = 8'hC9;
                    16'h7C4E: data_out = 8'hCA;
                    16'h7C4F: data_out = 8'hCB;
                    16'h7C50: data_out = 8'hCC;
                    16'h7C51: data_out = 8'hCD;
                    16'h7C52: data_out = 8'hCE;
                    16'h7C53: data_out = 8'hCF;
                    16'h7C54: data_out = 8'hD0;
                    16'h7C55: data_out = 8'hD1;
                    16'h7C56: data_out = 8'hD2;
                    16'h7C57: data_out = 8'hD3;
                    16'h7C58: data_out = 8'hD4;
                    16'h7C59: data_out = 8'hD5;
                    16'h7C5A: data_out = 8'hD6;
                    16'h7C5B: data_out = 8'hD7;
                    16'h7C5C: data_out = 8'hD8;
                    16'h7C5D: data_out = 8'hD9;
                    16'h7C5E: data_out = 8'hDA;
                    16'h7C5F: data_out = 8'hDB;
                    16'h7C60: data_out = 8'hDC;
                    16'h7C61: data_out = 8'hDD;
                    16'h7C62: data_out = 8'hDE;
                    16'h7C63: data_out = 8'hDF;
                    16'h7C64: data_out = 8'hE0;
                    16'h7C65: data_out = 8'hE1;
                    16'h7C66: data_out = 8'hE2;
                    16'h7C67: data_out = 8'hE3;
                    16'h7C68: data_out = 8'hE4;
                    16'h7C69: data_out = 8'hE5;
                    16'h7C6A: data_out = 8'hE6;
                    16'h7C6B: data_out = 8'hE7;
                    16'h7C6C: data_out = 8'hE8;
                    16'h7C6D: data_out = 8'hE9;
                    16'h7C6E: data_out = 8'hEA;
                    16'h7C6F: data_out = 8'hEB;
                    16'h7C70: data_out = 8'hEC;
                    16'h7C71: data_out = 8'hED;
                    16'h7C72: data_out = 8'hEE;
                    16'h7C73: data_out = 8'hEF;
                    16'h7C74: data_out = 8'hF0;
                    16'h7C75: data_out = 8'hF1;
                    16'h7C76: data_out = 8'hF2;
                    16'h7C77: data_out = 8'hF3;
                    16'h7C78: data_out = 8'hF4;
                    16'h7C79: data_out = 8'hF5;
                    16'h7C7A: data_out = 8'hF6;
                    16'h7C7B: data_out = 8'hF7;
                    16'h7C7C: data_out = 8'hF8;
                    16'h7C7D: data_out = 8'hF9;
                    16'h7C7E: data_out = 8'hFA;
                    16'h7C7F: data_out = 8'hFB;
                    16'h7C80: data_out = 8'h7C;
                    16'h7C81: data_out = 8'h7B;
                    16'h7C82: data_out = 8'h7A;
                    16'h7C83: data_out = 8'h79;
                    16'h7C84: data_out = 8'h78;
                    16'h7C85: data_out = 8'h77;
                    16'h7C86: data_out = 8'h76;
                    16'h7C87: data_out = 8'h75;
                    16'h7C88: data_out = 8'h74;
                    16'h7C89: data_out = 8'h73;
                    16'h7C8A: data_out = 8'h72;
                    16'h7C8B: data_out = 8'h71;
                    16'h7C8C: data_out = 8'h70;
                    16'h7C8D: data_out = 8'h6F;
                    16'h7C8E: data_out = 8'h6E;
                    16'h7C8F: data_out = 8'h6D;
                    16'h7C90: data_out = 8'h6C;
                    16'h7C91: data_out = 8'h6B;
                    16'h7C92: data_out = 8'h6A;
                    16'h7C93: data_out = 8'h69;
                    16'h7C94: data_out = 8'h68;
                    16'h7C95: data_out = 8'h67;
                    16'h7C96: data_out = 8'h66;
                    16'h7C97: data_out = 8'h65;
                    16'h7C98: data_out = 8'h64;
                    16'h7C99: data_out = 8'h63;
                    16'h7C9A: data_out = 8'h62;
                    16'h7C9B: data_out = 8'h61;
                    16'h7C9C: data_out = 8'h60;
                    16'h7C9D: data_out = 8'h5F;
                    16'h7C9E: data_out = 8'h5E;
                    16'h7C9F: data_out = 8'h5D;
                    16'h7CA0: data_out = 8'h5C;
                    16'h7CA1: data_out = 8'h5B;
                    16'h7CA2: data_out = 8'h5A;
                    16'h7CA3: data_out = 8'h59;
                    16'h7CA4: data_out = 8'h58;
                    16'h7CA5: data_out = 8'h57;
                    16'h7CA6: data_out = 8'h56;
                    16'h7CA7: data_out = 8'h55;
                    16'h7CA8: data_out = 8'h54;
                    16'h7CA9: data_out = 8'h53;
                    16'h7CAA: data_out = 8'h52;
                    16'h7CAB: data_out = 8'h51;
                    16'h7CAC: data_out = 8'h50;
                    16'h7CAD: data_out = 8'h4F;
                    16'h7CAE: data_out = 8'h4E;
                    16'h7CAF: data_out = 8'h4D;
                    16'h7CB0: data_out = 8'h4C;
                    16'h7CB1: data_out = 8'h4B;
                    16'h7CB2: data_out = 8'h4A;
                    16'h7CB3: data_out = 8'h49;
                    16'h7CB4: data_out = 8'h48;
                    16'h7CB5: data_out = 8'h47;
                    16'h7CB6: data_out = 8'h46;
                    16'h7CB7: data_out = 8'h45;
                    16'h7CB8: data_out = 8'h44;
                    16'h7CB9: data_out = 8'h43;
                    16'h7CBA: data_out = 8'h42;
                    16'h7CBB: data_out = 8'h41;
                    16'h7CBC: data_out = 8'h40;
                    16'h7CBD: data_out = 8'h3F;
                    16'h7CBE: data_out = 8'h3E;
                    16'h7CBF: data_out = 8'h3D;
                    16'h7CC0: data_out = 8'h3C;
                    16'h7CC1: data_out = 8'h3B;
                    16'h7CC2: data_out = 8'h3A;
                    16'h7CC3: data_out = 8'h39;
                    16'h7CC4: data_out = 8'h38;
                    16'h7CC5: data_out = 8'h37;
                    16'h7CC6: data_out = 8'h36;
                    16'h7CC7: data_out = 8'h35;
                    16'h7CC8: data_out = 8'h34;
                    16'h7CC9: data_out = 8'h33;
                    16'h7CCA: data_out = 8'h32;
                    16'h7CCB: data_out = 8'h31;
                    16'h7CCC: data_out = 8'h30;
                    16'h7CCD: data_out = 8'h2F;
                    16'h7CCE: data_out = 8'h2E;
                    16'h7CCF: data_out = 8'h2D;
                    16'h7CD0: data_out = 8'h2C;
                    16'h7CD1: data_out = 8'h2B;
                    16'h7CD2: data_out = 8'h2A;
                    16'h7CD3: data_out = 8'h29;
                    16'h7CD4: data_out = 8'h28;
                    16'h7CD5: data_out = 8'h27;
                    16'h7CD6: data_out = 8'h26;
                    16'h7CD7: data_out = 8'h25;
                    16'h7CD8: data_out = 8'h24;
                    16'h7CD9: data_out = 8'h23;
                    16'h7CDA: data_out = 8'h22;
                    16'h7CDB: data_out = 8'h21;
                    16'h7CDC: data_out = 8'h20;
                    16'h7CDD: data_out = 8'h1F;
                    16'h7CDE: data_out = 8'h1E;
                    16'h7CDF: data_out = 8'h1D;
                    16'h7CE0: data_out = 8'h1C;
                    16'h7CE1: data_out = 8'h1B;
                    16'h7CE2: data_out = 8'h1A;
                    16'h7CE3: data_out = 8'h19;
                    16'h7CE4: data_out = 8'h18;
                    16'h7CE5: data_out = 8'h17;
                    16'h7CE6: data_out = 8'h16;
                    16'h7CE7: data_out = 8'h15;
                    16'h7CE8: data_out = 8'h14;
                    16'h7CE9: data_out = 8'h13;
                    16'h7CEA: data_out = 8'h12;
                    16'h7CEB: data_out = 8'h11;
                    16'h7CEC: data_out = 8'h10;
                    16'h7CED: data_out = 8'hF;
                    16'h7CEE: data_out = 8'hE;
                    16'h7CEF: data_out = 8'hD;
                    16'h7CF0: data_out = 8'hC;
                    16'h7CF1: data_out = 8'hB;
                    16'h7CF2: data_out = 8'hA;
                    16'h7CF3: data_out = 8'h9;
                    16'h7CF4: data_out = 8'h8;
                    16'h7CF5: data_out = 8'h7;
                    16'h7CF6: data_out = 8'h6;
                    16'h7CF7: data_out = 8'h5;
                    16'h7CF8: data_out = 8'h4;
                    16'h7CF9: data_out = 8'h3;
                    16'h7CFA: data_out = 8'h2;
                    16'h7CFB: data_out = 8'h1;
                    16'h7CFC: data_out = 8'h0;
                    16'h7CFD: data_out = 8'h81;
                    16'h7CFE: data_out = 8'h82;
                    16'h7CFF: data_out = 8'h83;
                    16'h7D00: data_out = 8'h7D;
                    16'h7D01: data_out = 8'h7E;
                    16'h7D02: data_out = 8'h7F;
                    16'h7D03: data_out = 8'h80;
                    16'h7D04: data_out = 8'h81;
                    16'h7D05: data_out = 8'h82;
                    16'h7D06: data_out = 8'h83;
                    16'h7D07: data_out = 8'h84;
                    16'h7D08: data_out = 8'h85;
                    16'h7D09: data_out = 8'h86;
                    16'h7D0A: data_out = 8'h87;
                    16'h7D0B: data_out = 8'h88;
                    16'h7D0C: data_out = 8'h89;
                    16'h7D0D: data_out = 8'h8A;
                    16'h7D0E: data_out = 8'h8B;
                    16'h7D0F: data_out = 8'h8C;
                    16'h7D10: data_out = 8'h8D;
                    16'h7D11: data_out = 8'h8E;
                    16'h7D12: data_out = 8'h8F;
                    16'h7D13: data_out = 8'h90;
                    16'h7D14: data_out = 8'h91;
                    16'h7D15: data_out = 8'h92;
                    16'h7D16: data_out = 8'h93;
                    16'h7D17: data_out = 8'h94;
                    16'h7D18: data_out = 8'h95;
                    16'h7D19: data_out = 8'h96;
                    16'h7D1A: data_out = 8'h97;
                    16'h7D1B: data_out = 8'h98;
                    16'h7D1C: data_out = 8'h99;
                    16'h7D1D: data_out = 8'h9A;
                    16'h7D1E: data_out = 8'h9B;
                    16'h7D1F: data_out = 8'h9C;
                    16'h7D20: data_out = 8'h9D;
                    16'h7D21: data_out = 8'h9E;
                    16'h7D22: data_out = 8'h9F;
                    16'h7D23: data_out = 8'hA0;
                    16'h7D24: data_out = 8'hA1;
                    16'h7D25: data_out = 8'hA2;
                    16'h7D26: data_out = 8'hA3;
                    16'h7D27: data_out = 8'hA4;
                    16'h7D28: data_out = 8'hA5;
                    16'h7D29: data_out = 8'hA6;
                    16'h7D2A: data_out = 8'hA7;
                    16'h7D2B: data_out = 8'hA8;
                    16'h7D2C: data_out = 8'hA9;
                    16'h7D2D: data_out = 8'hAA;
                    16'h7D2E: data_out = 8'hAB;
                    16'h7D2F: data_out = 8'hAC;
                    16'h7D30: data_out = 8'hAD;
                    16'h7D31: data_out = 8'hAE;
                    16'h7D32: data_out = 8'hAF;
                    16'h7D33: data_out = 8'hB0;
                    16'h7D34: data_out = 8'hB1;
                    16'h7D35: data_out = 8'hB2;
                    16'h7D36: data_out = 8'hB3;
                    16'h7D37: data_out = 8'hB4;
                    16'h7D38: data_out = 8'hB5;
                    16'h7D39: data_out = 8'hB6;
                    16'h7D3A: data_out = 8'hB7;
                    16'h7D3B: data_out = 8'hB8;
                    16'h7D3C: data_out = 8'hB9;
                    16'h7D3D: data_out = 8'hBA;
                    16'h7D3E: data_out = 8'hBB;
                    16'h7D3F: data_out = 8'hBC;
                    16'h7D40: data_out = 8'hBD;
                    16'h7D41: data_out = 8'hBE;
                    16'h7D42: data_out = 8'hBF;
                    16'h7D43: data_out = 8'hC0;
                    16'h7D44: data_out = 8'hC1;
                    16'h7D45: data_out = 8'hC2;
                    16'h7D46: data_out = 8'hC3;
                    16'h7D47: data_out = 8'hC4;
                    16'h7D48: data_out = 8'hC5;
                    16'h7D49: data_out = 8'hC6;
                    16'h7D4A: data_out = 8'hC7;
                    16'h7D4B: data_out = 8'hC8;
                    16'h7D4C: data_out = 8'hC9;
                    16'h7D4D: data_out = 8'hCA;
                    16'h7D4E: data_out = 8'hCB;
                    16'h7D4F: data_out = 8'hCC;
                    16'h7D50: data_out = 8'hCD;
                    16'h7D51: data_out = 8'hCE;
                    16'h7D52: data_out = 8'hCF;
                    16'h7D53: data_out = 8'hD0;
                    16'h7D54: data_out = 8'hD1;
                    16'h7D55: data_out = 8'hD2;
                    16'h7D56: data_out = 8'hD3;
                    16'h7D57: data_out = 8'hD4;
                    16'h7D58: data_out = 8'hD5;
                    16'h7D59: data_out = 8'hD6;
                    16'h7D5A: data_out = 8'hD7;
                    16'h7D5B: data_out = 8'hD8;
                    16'h7D5C: data_out = 8'hD9;
                    16'h7D5D: data_out = 8'hDA;
                    16'h7D5E: data_out = 8'hDB;
                    16'h7D5F: data_out = 8'hDC;
                    16'h7D60: data_out = 8'hDD;
                    16'h7D61: data_out = 8'hDE;
                    16'h7D62: data_out = 8'hDF;
                    16'h7D63: data_out = 8'hE0;
                    16'h7D64: data_out = 8'hE1;
                    16'h7D65: data_out = 8'hE2;
                    16'h7D66: data_out = 8'hE3;
                    16'h7D67: data_out = 8'hE4;
                    16'h7D68: data_out = 8'hE5;
                    16'h7D69: data_out = 8'hE6;
                    16'h7D6A: data_out = 8'hE7;
                    16'h7D6B: data_out = 8'hE8;
                    16'h7D6C: data_out = 8'hE9;
                    16'h7D6D: data_out = 8'hEA;
                    16'h7D6E: data_out = 8'hEB;
                    16'h7D6F: data_out = 8'hEC;
                    16'h7D70: data_out = 8'hED;
                    16'h7D71: data_out = 8'hEE;
                    16'h7D72: data_out = 8'hEF;
                    16'h7D73: data_out = 8'hF0;
                    16'h7D74: data_out = 8'hF1;
                    16'h7D75: data_out = 8'hF2;
                    16'h7D76: data_out = 8'hF3;
                    16'h7D77: data_out = 8'hF4;
                    16'h7D78: data_out = 8'hF5;
                    16'h7D79: data_out = 8'hF6;
                    16'h7D7A: data_out = 8'hF7;
                    16'h7D7B: data_out = 8'hF8;
                    16'h7D7C: data_out = 8'hF9;
                    16'h7D7D: data_out = 8'hFA;
                    16'h7D7E: data_out = 8'hFB;
                    16'h7D7F: data_out = 8'hFC;
                    16'h7D80: data_out = 8'h7D;
                    16'h7D81: data_out = 8'h7C;
                    16'h7D82: data_out = 8'h7B;
                    16'h7D83: data_out = 8'h7A;
                    16'h7D84: data_out = 8'h79;
                    16'h7D85: data_out = 8'h78;
                    16'h7D86: data_out = 8'h77;
                    16'h7D87: data_out = 8'h76;
                    16'h7D88: data_out = 8'h75;
                    16'h7D89: data_out = 8'h74;
                    16'h7D8A: data_out = 8'h73;
                    16'h7D8B: data_out = 8'h72;
                    16'h7D8C: data_out = 8'h71;
                    16'h7D8D: data_out = 8'h70;
                    16'h7D8E: data_out = 8'h6F;
                    16'h7D8F: data_out = 8'h6E;
                    16'h7D90: data_out = 8'h6D;
                    16'h7D91: data_out = 8'h6C;
                    16'h7D92: data_out = 8'h6B;
                    16'h7D93: data_out = 8'h6A;
                    16'h7D94: data_out = 8'h69;
                    16'h7D95: data_out = 8'h68;
                    16'h7D96: data_out = 8'h67;
                    16'h7D97: data_out = 8'h66;
                    16'h7D98: data_out = 8'h65;
                    16'h7D99: data_out = 8'h64;
                    16'h7D9A: data_out = 8'h63;
                    16'h7D9B: data_out = 8'h62;
                    16'h7D9C: data_out = 8'h61;
                    16'h7D9D: data_out = 8'h60;
                    16'h7D9E: data_out = 8'h5F;
                    16'h7D9F: data_out = 8'h5E;
                    16'h7DA0: data_out = 8'h5D;
                    16'h7DA1: data_out = 8'h5C;
                    16'h7DA2: data_out = 8'h5B;
                    16'h7DA3: data_out = 8'h5A;
                    16'h7DA4: data_out = 8'h59;
                    16'h7DA5: data_out = 8'h58;
                    16'h7DA6: data_out = 8'h57;
                    16'h7DA7: data_out = 8'h56;
                    16'h7DA8: data_out = 8'h55;
                    16'h7DA9: data_out = 8'h54;
                    16'h7DAA: data_out = 8'h53;
                    16'h7DAB: data_out = 8'h52;
                    16'h7DAC: data_out = 8'h51;
                    16'h7DAD: data_out = 8'h50;
                    16'h7DAE: data_out = 8'h4F;
                    16'h7DAF: data_out = 8'h4E;
                    16'h7DB0: data_out = 8'h4D;
                    16'h7DB1: data_out = 8'h4C;
                    16'h7DB2: data_out = 8'h4B;
                    16'h7DB3: data_out = 8'h4A;
                    16'h7DB4: data_out = 8'h49;
                    16'h7DB5: data_out = 8'h48;
                    16'h7DB6: data_out = 8'h47;
                    16'h7DB7: data_out = 8'h46;
                    16'h7DB8: data_out = 8'h45;
                    16'h7DB9: data_out = 8'h44;
                    16'h7DBA: data_out = 8'h43;
                    16'h7DBB: data_out = 8'h42;
                    16'h7DBC: data_out = 8'h41;
                    16'h7DBD: data_out = 8'h40;
                    16'h7DBE: data_out = 8'h3F;
                    16'h7DBF: data_out = 8'h3E;
                    16'h7DC0: data_out = 8'h3D;
                    16'h7DC1: data_out = 8'h3C;
                    16'h7DC2: data_out = 8'h3B;
                    16'h7DC3: data_out = 8'h3A;
                    16'h7DC4: data_out = 8'h39;
                    16'h7DC5: data_out = 8'h38;
                    16'h7DC6: data_out = 8'h37;
                    16'h7DC7: data_out = 8'h36;
                    16'h7DC8: data_out = 8'h35;
                    16'h7DC9: data_out = 8'h34;
                    16'h7DCA: data_out = 8'h33;
                    16'h7DCB: data_out = 8'h32;
                    16'h7DCC: data_out = 8'h31;
                    16'h7DCD: data_out = 8'h30;
                    16'h7DCE: data_out = 8'h2F;
                    16'h7DCF: data_out = 8'h2E;
                    16'h7DD0: data_out = 8'h2D;
                    16'h7DD1: data_out = 8'h2C;
                    16'h7DD2: data_out = 8'h2B;
                    16'h7DD3: data_out = 8'h2A;
                    16'h7DD4: data_out = 8'h29;
                    16'h7DD5: data_out = 8'h28;
                    16'h7DD6: data_out = 8'h27;
                    16'h7DD7: data_out = 8'h26;
                    16'h7DD8: data_out = 8'h25;
                    16'h7DD9: data_out = 8'h24;
                    16'h7DDA: data_out = 8'h23;
                    16'h7DDB: data_out = 8'h22;
                    16'h7DDC: data_out = 8'h21;
                    16'h7DDD: data_out = 8'h20;
                    16'h7DDE: data_out = 8'h1F;
                    16'h7DDF: data_out = 8'h1E;
                    16'h7DE0: data_out = 8'h1D;
                    16'h7DE1: data_out = 8'h1C;
                    16'h7DE2: data_out = 8'h1B;
                    16'h7DE3: data_out = 8'h1A;
                    16'h7DE4: data_out = 8'h19;
                    16'h7DE5: data_out = 8'h18;
                    16'h7DE6: data_out = 8'h17;
                    16'h7DE7: data_out = 8'h16;
                    16'h7DE8: data_out = 8'h15;
                    16'h7DE9: data_out = 8'h14;
                    16'h7DEA: data_out = 8'h13;
                    16'h7DEB: data_out = 8'h12;
                    16'h7DEC: data_out = 8'h11;
                    16'h7DED: data_out = 8'h10;
                    16'h7DEE: data_out = 8'hF;
                    16'h7DEF: data_out = 8'hE;
                    16'h7DF0: data_out = 8'hD;
                    16'h7DF1: data_out = 8'hC;
                    16'h7DF2: data_out = 8'hB;
                    16'h7DF3: data_out = 8'hA;
                    16'h7DF4: data_out = 8'h9;
                    16'h7DF5: data_out = 8'h8;
                    16'h7DF6: data_out = 8'h7;
                    16'h7DF7: data_out = 8'h6;
                    16'h7DF8: data_out = 8'h5;
                    16'h7DF9: data_out = 8'h4;
                    16'h7DFA: data_out = 8'h3;
                    16'h7DFB: data_out = 8'h2;
                    16'h7DFC: data_out = 8'h1;
                    16'h7DFD: data_out = 8'h0;
                    16'h7DFE: data_out = 8'h81;
                    16'h7DFF: data_out = 8'h82;
                    16'h7E00: data_out = 8'h7E;
                    16'h7E01: data_out = 8'h7F;
                    16'h7E02: data_out = 8'h80;
                    16'h7E03: data_out = 8'h81;
                    16'h7E04: data_out = 8'h82;
                    16'h7E05: data_out = 8'h83;
                    16'h7E06: data_out = 8'h84;
                    16'h7E07: data_out = 8'h85;
                    16'h7E08: data_out = 8'h86;
                    16'h7E09: data_out = 8'h87;
                    16'h7E0A: data_out = 8'h88;
                    16'h7E0B: data_out = 8'h89;
                    16'h7E0C: data_out = 8'h8A;
                    16'h7E0D: data_out = 8'h8B;
                    16'h7E0E: data_out = 8'h8C;
                    16'h7E0F: data_out = 8'h8D;
                    16'h7E10: data_out = 8'h8E;
                    16'h7E11: data_out = 8'h8F;
                    16'h7E12: data_out = 8'h90;
                    16'h7E13: data_out = 8'h91;
                    16'h7E14: data_out = 8'h92;
                    16'h7E15: data_out = 8'h93;
                    16'h7E16: data_out = 8'h94;
                    16'h7E17: data_out = 8'h95;
                    16'h7E18: data_out = 8'h96;
                    16'h7E19: data_out = 8'h97;
                    16'h7E1A: data_out = 8'h98;
                    16'h7E1B: data_out = 8'h99;
                    16'h7E1C: data_out = 8'h9A;
                    16'h7E1D: data_out = 8'h9B;
                    16'h7E1E: data_out = 8'h9C;
                    16'h7E1F: data_out = 8'h9D;
                    16'h7E20: data_out = 8'h9E;
                    16'h7E21: data_out = 8'h9F;
                    16'h7E22: data_out = 8'hA0;
                    16'h7E23: data_out = 8'hA1;
                    16'h7E24: data_out = 8'hA2;
                    16'h7E25: data_out = 8'hA3;
                    16'h7E26: data_out = 8'hA4;
                    16'h7E27: data_out = 8'hA5;
                    16'h7E28: data_out = 8'hA6;
                    16'h7E29: data_out = 8'hA7;
                    16'h7E2A: data_out = 8'hA8;
                    16'h7E2B: data_out = 8'hA9;
                    16'h7E2C: data_out = 8'hAA;
                    16'h7E2D: data_out = 8'hAB;
                    16'h7E2E: data_out = 8'hAC;
                    16'h7E2F: data_out = 8'hAD;
                    16'h7E30: data_out = 8'hAE;
                    16'h7E31: data_out = 8'hAF;
                    16'h7E32: data_out = 8'hB0;
                    16'h7E33: data_out = 8'hB1;
                    16'h7E34: data_out = 8'hB2;
                    16'h7E35: data_out = 8'hB3;
                    16'h7E36: data_out = 8'hB4;
                    16'h7E37: data_out = 8'hB5;
                    16'h7E38: data_out = 8'hB6;
                    16'h7E39: data_out = 8'hB7;
                    16'h7E3A: data_out = 8'hB8;
                    16'h7E3B: data_out = 8'hB9;
                    16'h7E3C: data_out = 8'hBA;
                    16'h7E3D: data_out = 8'hBB;
                    16'h7E3E: data_out = 8'hBC;
                    16'h7E3F: data_out = 8'hBD;
                    16'h7E40: data_out = 8'hBE;
                    16'h7E41: data_out = 8'hBF;
                    16'h7E42: data_out = 8'hC0;
                    16'h7E43: data_out = 8'hC1;
                    16'h7E44: data_out = 8'hC2;
                    16'h7E45: data_out = 8'hC3;
                    16'h7E46: data_out = 8'hC4;
                    16'h7E47: data_out = 8'hC5;
                    16'h7E48: data_out = 8'hC6;
                    16'h7E49: data_out = 8'hC7;
                    16'h7E4A: data_out = 8'hC8;
                    16'h7E4B: data_out = 8'hC9;
                    16'h7E4C: data_out = 8'hCA;
                    16'h7E4D: data_out = 8'hCB;
                    16'h7E4E: data_out = 8'hCC;
                    16'h7E4F: data_out = 8'hCD;
                    16'h7E50: data_out = 8'hCE;
                    16'h7E51: data_out = 8'hCF;
                    16'h7E52: data_out = 8'hD0;
                    16'h7E53: data_out = 8'hD1;
                    16'h7E54: data_out = 8'hD2;
                    16'h7E55: data_out = 8'hD3;
                    16'h7E56: data_out = 8'hD4;
                    16'h7E57: data_out = 8'hD5;
                    16'h7E58: data_out = 8'hD6;
                    16'h7E59: data_out = 8'hD7;
                    16'h7E5A: data_out = 8'hD8;
                    16'h7E5B: data_out = 8'hD9;
                    16'h7E5C: data_out = 8'hDA;
                    16'h7E5D: data_out = 8'hDB;
                    16'h7E5E: data_out = 8'hDC;
                    16'h7E5F: data_out = 8'hDD;
                    16'h7E60: data_out = 8'hDE;
                    16'h7E61: data_out = 8'hDF;
                    16'h7E62: data_out = 8'hE0;
                    16'h7E63: data_out = 8'hE1;
                    16'h7E64: data_out = 8'hE2;
                    16'h7E65: data_out = 8'hE3;
                    16'h7E66: data_out = 8'hE4;
                    16'h7E67: data_out = 8'hE5;
                    16'h7E68: data_out = 8'hE6;
                    16'h7E69: data_out = 8'hE7;
                    16'h7E6A: data_out = 8'hE8;
                    16'h7E6B: data_out = 8'hE9;
                    16'h7E6C: data_out = 8'hEA;
                    16'h7E6D: data_out = 8'hEB;
                    16'h7E6E: data_out = 8'hEC;
                    16'h7E6F: data_out = 8'hED;
                    16'h7E70: data_out = 8'hEE;
                    16'h7E71: data_out = 8'hEF;
                    16'h7E72: data_out = 8'hF0;
                    16'h7E73: data_out = 8'hF1;
                    16'h7E74: data_out = 8'hF2;
                    16'h7E75: data_out = 8'hF3;
                    16'h7E76: data_out = 8'hF4;
                    16'h7E77: data_out = 8'hF5;
                    16'h7E78: data_out = 8'hF6;
                    16'h7E79: data_out = 8'hF7;
                    16'h7E7A: data_out = 8'hF8;
                    16'h7E7B: data_out = 8'hF9;
                    16'h7E7C: data_out = 8'hFA;
                    16'h7E7D: data_out = 8'hFB;
                    16'h7E7E: data_out = 8'hFC;
                    16'h7E7F: data_out = 8'hFD;
                    16'h7E80: data_out = 8'h7E;
                    16'h7E81: data_out = 8'h7D;
                    16'h7E82: data_out = 8'h7C;
                    16'h7E83: data_out = 8'h7B;
                    16'h7E84: data_out = 8'h7A;
                    16'h7E85: data_out = 8'h79;
                    16'h7E86: data_out = 8'h78;
                    16'h7E87: data_out = 8'h77;
                    16'h7E88: data_out = 8'h76;
                    16'h7E89: data_out = 8'h75;
                    16'h7E8A: data_out = 8'h74;
                    16'h7E8B: data_out = 8'h73;
                    16'h7E8C: data_out = 8'h72;
                    16'h7E8D: data_out = 8'h71;
                    16'h7E8E: data_out = 8'h70;
                    16'h7E8F: data_out = 8'h6F;
                    16'h7E90: data_out = 8'h6E;
                    16'h7E91: data_out = 8'h6D;
                    16'h7E92: data_out = 8'h6C;
                    16'h7E93: data_out = 8'h6B;
                    16'h7E94: data_out = 8'h6A;
                    16'h7E95: data_out = 8'h69;
                    16'h7E96: data_out = 8'h68;
                    16'h7E97: data_out = 8'h67;
                    16'h7E98: data_out = 8'h66;
                    16'h7E99: data_out = 8'h65;
                    16'h7E9A: data_out = 8'h64;
                    16'h7E9B: data_out = 8'h63;
                    16'h7E9C: data_out = 8'h62;
                    16'h7E9D: data_out = 8'h61;
                    16'h7E9E: data_out = 8'h60;
                    16'h7E9F: data_out = 8'h5F;
                    16'h7EA0: data_out = 8'h5E;
                    16'h7EA1: data_out = 8'h5D;
                    16'h7EA2: data_out = 8'h5C;
                    16'h7EA3: data_out = 8'h5B;
                    16'h7EA4: data_out = 8'h5A;
                    16'h7EA5: data_out = 8'h59;
                    16'h7EA6: data_out = 8'h58;
                    16'h7EA7: data_out = 8'h57;
                    16'h7EA8: data_out = 8'h56;
                    16'h7EA9: data_out = 8'h55;
                    16'h7EAA: data_out = 8'h54;
                    16'h7EAB: data_out = 8'h53;
                    16'h7EAC: data_out = 8'h52;
                    16'h7EAD: data_out = 8'h51;
                    16'h7EAE: data_out = 8'h50;
                    16'h7EAF: data_out = 8'h4F;
                    16'h7EB0: data_out = 8'h4E;
                    16'h7EB1: data_out = 8'h4D;
                    16'h7EB2: data_out = 8'h4C;
                    16'h7EB3: data_out = 8'h4B;
                    16'h7EB4: data_out = 8'h4A;
                    16'h7EB5: data_out = 8'h49;
                    16'h7EB6: data_out = 8'h48;
                    16'h7EB7: data_out = 8'h47;
                    16'h7EB8: data_out = 8'h46;
                    16'h7EB9: data_out = 8'h45;
                    16'h7EBA: data_out = 8'h44;
                    16'h7EBB: data_out = 8'h43;
                    16'h7EBC: data_out = 8'h42;
                    16'h7EBD: data_out = 8'h41;
                    16'h7EBE: data_out = 8'h40;
                    16'h7EBF: data_out = 8'h3F;
                    16'h7EC0: data_out = 8'h3E;
                    16'h7EC1: data_out = 8'h3D;
                    16'h7EC2: data_out = 8'h3C;
                    16'h7EC3: data_out = 8'h3B;
                    16'h7EC4: data_out = 8'h3A;
                    16'h7EC5: data_out = 8'h39;
                    16'h7EC6: data_out = 8'h38;
                    16'h7EC7: data_out = 8'h37;
                    16'h7EC8: data_out = 8'h36;
                    16'h7EC9: data_out = 8'h35;
                    16'h7ECA: data_out = 8'h34;
                    16'h7ECB: data_out = 8'h33;
                    16'h7ECC: data_out = 8'h32;
                    16'h7ECD: data_out = 8'h31;
                    16'h7ECE: data_out = 8'h30;
                    16'h7ECF: data_out = 8'h2F;
                    16'h7ED0: data_out = 8'h2E;
                    16'h7ED1: data_out = 8'h2D;
                    16'h7ED2: data_out = 8'h2C;
                    16'h7ED3: data_out = 8'h2B;
                    16'h7ED4: data_out = 8'h2A;
                    16'h7ED5: data_out = 8'h29;
                    16'h7ED6: data_out = 8'h28;
                    16'h7ED7: data_out = 8'h27;
                    16'h7ED8: data_out = 8'h26;
                    16'h7ED9: data_out = 8'h25;
                    16'h7EDA: data_out = 8'h24;
                    16'h7EDB: data_out = 8'h23;
                    16'h7EDC: data_out = 8'h22;
                    16'h7EDD: data_out = 8'h21;
                    16'h7EDE: data_out = 8'h20;
                    16'h7EDF: data_out = 8'h1F;
                    16'h7EE0: data_out = 8'h1E;
                    16'h7EE1: data_out = 8'h1D;
                    16'h7EE2: data_out = 8'h1C;
                    16'h7EE3: data_out = 8'h1B;
                    16'h7EE4: data_out = 8'h1A;
                    16'h7EE5: data_out = 8'h19;
                    16'h7EE6: data_out = 8'h18;
                    16'h7EE7: data_out = 8'h17;
                    16'h7EE8: data_out = 8'h16;
                    16'h7EE9: data_out = 8'h15;
                    16'h7EEA: data_out = 8'h14;
                    16'h7EEB: data_out = 8'h13;
                    16'h7EEC: data_out = 8'h12;
                    16'h7EED: data_out = 8'h11;
                    16'h7EEE: data_out = 8'h10;
                    16'h7EEF: data_out = 8'hF;
                    16'h7EF0: data_out = 8'hE;
                    16'h7EF1: data_out = 8'hD;
                    16'h7EF2: data_out = 8'hC;
                    16'h7EF3: data_out = 8'hB;
                    16'h7EF4: data_out = 8'hA;
                    16'h7EF5: data_out = 8'h9;
                    16'h7EF6: data_out = 8'h8;
                    16'h7EF7: data_out = 8'h7;
                    16'h7EF8: data_out = 8'h6;
                    16'h7EF9: data_out = 8'h5;
                    16'h7EFA: data_out = 8'h4;
                    16'h7EFB: data_out = 8'h3;
                    16'h7EFC: data_out = 8'h2;
                    16'h7EFD: data_out = 8'h1;
                    16'h7EFE: data_out = 8'h0;
                    16'h7EFF: data_out = 8'h81;
                    16'h7F00: data_out = 8'h7F;
                    16'h7F01: data_out = 8'h80;
                    16'h7F02: data_out = 8'h81;
                    16'h7F03: data_out = 8'h82;
                    16'h7F04: data_out = 8'h83;
                    16'h7F05: data_out = 8'h84;
                    16'h7F06: data_out = 8'h85;
                    16'h7F07: data_out = 8'h86;
                    16'h7F08: data_out = 8'h87;
                    16'h7F09: data_out = 8'h88;
                    16'h7F0A: data_out = 8'h89;
                    16'h7F0B: data_out = 8'h8A;
                    16'h7F0C: data_out = 8'h8B;
                    16'h7F0D: data_out = 8'h8C;
                    16'h7F0E: data_out = 8'h8D;
                    16'h7F0F: data_out = 8'h8E;
                    16'h7F10: data_out = 8'h8F;
                    16'h7F11: data_out = 8'h90;
                    16'h7F12: data_out = 8'h91;
                    16'h7F13: data_out = 8'h92;
                    16'h7F14: data_out = 8'h93;
                    16'h7F15: data_out = 8'h94;
                    16'h7F16: data_out = 8'h95;
                    16'h7F17: data_out = 8'h96;
                    16'h7F18: data_out = 8'h97;
                    16'h7F19: data_out = 8'h98;
                    16'h7F1A: data_out = 8'h99;
                    16'h7F1B: data_out = 8'h9A;
                    16'h7F1C: data_out = 8'h9B;
                    16'h7F1D: data_out = 8'h9C;
                    16'h7F1E: data_out = 8'h9D;
                    16'h7F1F: data_out = 8'h9E;
                    16'h7F20: data_out = 8'h9F;
                    16'h7F21: data_out = 8'hA0;
                    16'h7F22: data_out = 8'hA1;
                    16'h7F23: data_out = 8'hA2;
                    16'h7F24: data_out = 8'hA3;
                    16'h7F25: data_out = 8'hA4;
                    16'h7F26: data_out = 8'hA5;
                    16'h7F27: data_out = 8'hA6;
                    16'h7F28: data_out = 8'hA7;
                    16'h7F29: data_out = 8'hA8;
                    16'h7F2A: data_out = 8'hA9;
                    16'h7F2B: data_out = 8'hAA;
                    16'h7F2C: data_out = 8'hAB;
                    16'h7F2D: data_out = 8'hAC;
                    16'h7F2E: data_out = 8'hAD;
                    16'h7F2F: data_out = 8'hAE;
                    16'h7F30: data_out = 8'hAF;
                    16'h7F31: data_out = 8'hB0;
                    16'h7F32: data_out = 8'hB1;
                    16'h7F33: data_out = 8'hB2;
                    16'h7F34: data_out = 8'hB3;
                    16'h7F35: data_out = 8'hB4;
                    16'h7F36: data_out = 8'hB5;
                    16'h7F37: data_out = 8'hB6;
                    16'h7F38: data_out = 8'hB7;
                    16'h7F39: data_out = 8'hB8;
                    16'h7F3A: data_out = 8'hB9;
                    16'h7F3B: data_out = 8'hBA;
                    16'h7F3C: data_out = 8'hBB;
                    16'h7F3D: data_out = 8'hBC;
                    16'h7F3E: data_out = 8'hBD;
                    16'h7F3F: data_out = 8'hBE;
                    16'h7F40: data_out = 8'hBF;
                    16'h7F41: data_out = 8'hC0;
                    16'h7F42: data_out = 8'hC1;
                    16'h7F43: data_out = 8'hC2;
                    16'h7F44: data_out = 8'hC3;
                    16'h7F45: data_out = 8'hC4;
                    16'h7F46: data_out = 8'hC5;
                    16'h7F47: data_out = 8'hC6;
                    16'h7F48: data_out = 8'hC7;
                    16'h7F49: data_out = 8'hC8;
                    16'h7F4A: data_out = 8'hC9;
                    16'h7F4B: data_out = 8'hCA;
                    16'h7F4C: data_out = 8'hCB;
                    16'h7F4D: data_out = 8'hCC;
                    16'h7F4E: data_out = 8'hCD;
                    16'h7F4F: data_out = 8'hCE;
                    16'h7F50: data_out = 8'hCF;
                    16'h7F51: data_out = 8'hD0;
                    16'h7F52: data_out = 8'hD1;
                    16'h7F53: data_out = 8'hD2;
                    16'h7F54: data_out = 8'hD3;
                    16'h7F55: data_out = 8'hD4;
                    16'h7F56: data_out = 8'hD5;
                    16'h7F57: data_out = 8'hD6;
                    16'h7F58: data_out = 8'hD7;
                    16'h7F59: data_out = 8'hD8;
                    16'h7F5A: data_out = 8'hD9;
                    16'h7F5B: data_out = 8'hDA;
                    16'h7F5C: data_out = 8'hDB;
                    16'h7F5D: data_out = 8'hDC;
                    16'h7F5E: data_out = 8'hDD;
                    16'h7F5F: data_out = 8'hDE;
                    16'h7F60: data_out = 8'hDF;
                    16'h7F61: data_out = 8'hE0;
                    16'h7F62: data_out = 8'hE1;
                    16'h7F63: data_out = 8'hE2;
                    16'h7F64: data_out = 8'hE3;
                    16'h7F65: data_out = 8'hE4;
                    16'h7F66: data_out = 8'hE5;
                    16'h7F67: data_out = 8'hE6;
                    16'h7F68: data_out = 8'hE7;
                    16'h7F69: data_out = 8'hE8;
                    16'h7F6A: data_out = 8'hE9;
                    16'h7F6B: data_out = 8'hEA;
                    16'h7F6C: data_out = 8'hEB;
                    16'h7F6D: data_out = 8'hEC;
                    16'h7F6E: data_out = 8'hED;
                    16'h7F6F: data_out = 8'hEE;
                    16'h7F70: data_out = 8'hEF;
                    16'h7F71: data_out = 8'hF0;
                    16'h7F72: data_out = 8'hF1;
                    16'h7F73: data_out = 8'hF2;
                    16'h7F74: data_out = 8'hF3;
                    16'h7F75: data_out = 8'hF4;
                    16'h7F76: data_out = 8'hF5;
                    16'h7F77: data_out = 8'hF6;
                    16'h7F78: data_out = 8'hF7;
                    16'h7F79: data_out = 8'hF8;
                    16'h7F7A: data_out = 8'hF9;
                    16'h7F7B: data_out = 8'hFA;
                    16'h7F7C: data_out = 8'hFB;
                    16'h7F7D: data_out = 8'hFC;
                    16'h7F7E: data_out = 8'hFD;
                    16'h7F7F: data_out = 8'hFE;
                    16'h7F80: data_out = 8'h7F;
                    16'h7F81: data_out = 8'h7E;
                    16'h7F82: data_out = 8'h7D;
                    16'h7F83: data_out = 8'h7C;
                    16'h7F84: data_out = 8'h7B;
                    16'h7F85: data_out = 8'h7A;
                    16'h7F86: data_out = 8'h79;
                    16'h7F87: data_out = 8'h78;
                    16'h7F88: data_out = 8'h77;
                    16'h7F89: data_out = 8'h76;
                    16'h7F8A: data_out = 8'h75;
                    16'h7F8B: data_out = 8'h74;
                    16'h7F8C: data_out = 8'h73;
                    16'h7F8D: data_out = 8'h72;
                    16'h7F8E: data_out = 8'h71;
                    16'h7F8F: data_out = 8'h70;
                    16'h7F90: data_out = 8'h6F;
                    16'h7F91: data_out = 8'h6E;
                    16'h7F92: data_out = 8'h6D;
                    16'h7F93: data_out = 8'h6C;
                    16'h7F94: data_out = 8'h6B;
                    16'h7F95: data_out = 8'h6A;
                    16'h7F96: data_out = 8'h69;
                    16'h7F97: data_out = 8'h68;
                    16'h7F98: data_out = 8'h67;
                    16'h7F99: data_out = 8'h66;
                    16'h7F9A: data_out = 8'h65;
                    16'h7F9B: data_out = 8'h64;
                    16'h7F9C: data_out = 8'h63;
                    16'h7F9D: data_out = 8'h62;
                    16'h7F9E: data_out = 8'h61;
                    16'h7F9F: data_out = 8'h60;
                    16'h7FA0: data_out = 8'h5F;
                    16'h7FA1: data_out = 8'h5E;
                    16'h7FA2: data_out = 8'h5D;
                    16'h7FA3: data_out = 8'h5C;
                    16'h7FA4: data_out = 8'h5B;
                    16'h7FA5: data_out = 8'h5A;
                    16'h7FA6: data_out = 8'h59;
                    16'h7FA7: data_out = 8'h58;
                    16'h7FA8: data_out = 8'h57;
                    16'h7FA9: data_out = 8'h56;
                    16'h7FAA: data_out = 8'h55;
                    16'h7FAB: data_out = 8'h54;
                    16'h7FAC: data_out = 8'h53;
                    16'h7FAD: data_out = 8'h52;
                    16'h7FAE: data_out = 8'h51;
                    16'h7FAF: data_out = 8'h50;
                    16'h7FB0: data_out = 8'h4F;
                    16'h7FB1: data_out = 8'h4E;
                    16'h7FB2: data_out = 8'h4D;
                    16'h7FB3: data_out = 8'h4C;
                    16'h7FB4: data_out = 8'h4B;
                    16'h7FB5: data_out = 8'h4A;
                    16'h7FB6: data_out = 8'h49;
                    16'h7FB7: data_out = 8'h48;
                    16'h7FB8: data_out = 8'h47;
                    16'h7FB9: data_out = 8'h46;
                    16'h7FBA: data_out = 8'h45;
                    16'h7FBB: data_out = 8'h44;
                    16'h7FBC: data_out = 8'h43;
                    16'h7FBD: data_out = 8'h42;
                    16'h7FBE: data_out = 8'h41;
                    16'h7FBF: data_out = 8'h40;
                    16'h7FC0: data_out = 8'h3F;
                    16'h7FC1: data_out = 8'h3E;
                    16'h7FC2: data_out = 8'h3D;
                    16'h7FC3: data_out = 8'h3C;
                    16'h7FC4: data_out = 8'h3B;
                    16'h7FC5: data_out = 8'h3A;
                    16'h7FC6: data_out = 8'h39;
                    16'h7FC7: data_out = 8'h38;
                    16'h7FC8: data_out = 8'h37;
                    16'h7FC9: data_out = 8'h36;
                    16'h7FCA: data_out = 8'h35;
                    16'h7FCB: data_out = 8'h34;
                    16'h7FCC: data_out = 8'h33;
                    16'h7FCD: data_out = 8'h32;
                    16'h7FCE: data_out = 8'h31;
                    16'h7FCF: data_out = 8'h30;
                    16'h7FD0: data_out = 8'h2F;
                    16'h7FD1: data_out = 8'h2E;
                    16'h7FD2: data_out = 8'h2D;
                    16'h7FD3: data_out = 8'h2C;
                    16'h7FD4: data_out = 8'h2B;
                    16'h7FD5: data_out = 8'h2A;
                    16'h7FD6: data_out = 8'h29;
                    16'h7FD7: data_out = 8'h28;
                    16'h7FD8: data_out = 8'h27;
                    16'h7FD9: data_out = 8'h26;
                    16'h7FDA: data_out = 8'h25;
                    16'h7FDB: data_out = 8'h24;
                    16'h7FDC: data_out = 8'h23;
                    16'h7FDD: data_out = 8'h22;
                    16'h7FDE: data_out = 8'h21;
                    16'h7FDF: data_out = 8'h20;
                    16'h7FE0: data_out = 8'h1F;
                    16'h7FE1: data_out = 8'h1E;
                    16'h7FE2: data_out = 8'h1D;
                    16'h7FE3: data_out = 8'h1C;
                    16'h7FE4: data_out = 8'h1B;
                    16'h7FE5: data_out = 8'h1A;
                    16'h7FE6: data_out = 8'h19;
                    16'h7FE7: data_out = 8'h18;
                    16'h7FE8: data_out = 8'h17;
                    16'h7FE9: data_out = 8'h16;
                    16'h7FEA: data_out = 8'h15;
                    16'h7FEB: data_out = 8'h14;
                    16'h7FEC: data_out = 8'h13;
                    16'h7FED: data_out = 8'h12;
                    16'h7FEE: data_out = 8'h11;
                    16'h7FEF: data_out = 8'h10;
                    16'h7FF0: data_out = 8'hF;
                    16'h7FF1: data_out = 8'hE;
                    16'h7FF2: data_out = 8'hD;
                    16'h7FF3: data_out = 8'hC;
                    16'h7FF4: data_out = 8'hB;
                    16'h7FF5: data_out = 8'hA;
                    16'h7FF6: data_out = 8'h9;
                    16'h7FF7: data_out = 8'h8;
                    16'h7FF8: data_out = 8'h7;
                    16'h7FF9: data_out = 8'h6;
                    16'h7FFA: data_out = 8'h5;
                    16'h7FFB: data_out = 8'h4;
                    16'h7FFC: data_out = 8'h3;
                    16'h7FFD: data_out = 8'h2;
                    16'h7FFE: data_out = 8'h1;
                    16'h7FFF: data_out = 8'h0;
                    16'h8000: data_out = 8'h0;
                    16'h8001: data_out = 8'h1;
                    16'h8002: data_out = 8'h2;
                    16'h8003: data_out = 8'h3;
                    16'h8004: data_out = 8'h4;
                    16'h8005: data_out = 8'h5;
                    16'h8006: data_out = 8'h6;
                    16'h8007: data_out = 8'h7;
                    16'h8008: data_out = 8'h8;
                    16'h8009: data_out = 8'h9;
                    16'h800A: data_out = 8'hA;
                    16'h800B: data_out = 8'hB;
                    16'h800C: data_out = 8'hC;
                    16'h800D: data_out = 8'hD;
                    16'h800E: data_out = 8'hE;
                    16'h800F: data_out = 8'hF;
                    16'h8010: data_out = 8'h10;
                    16'h8011: data_out = 8'h11;
                    16'h8012: data_out = 8'h12;
                    16'h8013: data_out = 8'h13;
                    16'h8014: data_out = 8'h14;
                    16'h8015: data_out = 8'h15;
                    16'h8016: data_out = 8'h16;
                    16'h8017: data_out = 8'h17;
                    16'h8018: data_out = 8'h18;
                    16'h8019: data_out = 8'h19;
                    16'h801A: data_out = 8'h1A;
                    16'h801B: data_out = 8'h1B;
                    16'h801C: data_out = 8'h1C;
                    16'h801D: data_out = 8'h1D;
                    16'h801E: data_out = 8'h1E;
                    16'h801F: data_out = 8'h1F;
                    16'h8020: data_out = 8'h20;
                    16'h8021: data_out = 8'h21;
                    16'h8022: data_out = 8'h22;
                    16'h8023: data_out = 8'h23;
                    16'h8024: data_out = 8'h24;
                    16'h8025: data_out = 8'h25;
                    16'h8026: data_out = 8'h26;
                    16'h8027: data_out = 8'h27;
                    16'h8028: data_out = 8'h28;
                    16'h8029: data_out = 8'h29;
                    16'h802A: data_out = 8'h2A;
                    16'h802B: data_out = 8'h2B;
                    16'h802C: data_out = 8'h2C;
                    16'h802D: data_out = 8'h2D;
                    16'h802E: data_out = 8'h2E;
                    16'h802F: data_out = 8'h2F;
                    16'h8030: data_out = 8'h30;
                    16'h8031: data_out = 8'h31;
                    16'h8032: data_out = 8'h32;
                    16'h8033: data_out = 8'h33;
                    16'h8034: data_out = 8'h34;
                    16'h8035: data_out = 8'h35;
                    16'h8036: data_out = 8'h36;
                    16'h8037: data_out = 8'h37;
                    16'h8038: data_out = 8'h38;
                    16'h8039: data_out = 8'h39;
                    16'h803A: data_out = 8'h3A;
                    16'h803B: data_out = 8'h3B;
                    16'h803C: data_out = 8'h3C;
                    16'h803D: data_out = 8'h3D;
                    16'h803E: data_out = 8'h3E;
                    16'h803F: data_out = 8'h3F;
                    16'h8040: data_out = 8'h40;
                    16'h8041: data_out = 8'h41;
                    16'h8042: data_out = 8'h42;
                    16'h8043: data_out = 8'h43;
                    16'h8044: data_out = 8'h44;
                    16'h8045: data_out = 8'h45;
                    16'h8046: data_out = 8'h46;
                    16'h8047: data_out = 8'h47;
                    16'h8048: data_out = 8'h48;
                    16'h8049: data_out = 8'h49;
                    16'h804A: data_out = 8'h4A;
                    16'h804B: data_out = 8'h4B;
                    16'h804C: data_out = 8'h4C;
                    16'h804D: data_out = 8'h4D;
                    16'h804E: data_out = 8'h4E;
                    16'h804F: data_out = 8'h4F;
                    16'h8050: data_out = 8'h50;
                    16'h8051: data_out = 8'h51;
                    16'h8052: data_out = 8'h52;
                    16'h8053: data_out = 8'h53;
                    16'h8054: data_out = 8'h54;
                    16'h8055: data_out = 8'h55;
                    16'h8056: data_out = 8'h56;
                    16'h8057: data_out = 8'h57;
                    16'h8058: data_out = 8'h58;
                    16'h8059: data_out = 8'h59;
                    16'h805A: data_out = 8'h5A;
                    16'h805B: data_out = 8'h5B;
                    16'h805C: data_out = 8'h5C;
                    16'h805D: data_out = 8'h5D;
                    16'h805E: data_out = 8'h5E;
                    16'h805F: data_out = 8'h5F;
                    16'h8060: data_out = 8'h60;
                    16'h8061: data_out = 8'h61;
                    16'h8062: data_out = 8'h62;
                    16'h8063: data_out = 8'h63;
                    16'h8064: data_out = 8'h64;
                    16'h8065: data_out = 8'h65;
                    16'h8066: data_out = 8'h66;
                    16'h8067: data_out = 8'h67;
                    16'h8068: data_out = 8'h68;
                    16'h8069: data_out = 8'h69;
                    16'h806A: data_out = 8'h6A;
                    16'h806B: data_out = 8'h6B;
                    16'h806C: data_out = 8'h6C;
                    16'h806D: data_out = 8'h6D;
                    16'h806E: data_out = 8'h6E;
                    16'h806F: data_out = 8'h6F;
                    16'h8070: data_out = 8'h70;
                    16'h8071: data_out = 8'h71;
                    16'h8072: data_out = 8'h72;
                    16'h8073: data_out = 8'h73;
                    16'h8074: data_out = 8'h74;
                    16'h8075: data_out = 8'h75;
                    16'h8076: data_out = 8'h76;
                    16'h8077: data_out = 8'h77;
                    16'h8078: data_out = 8'h78;
                    16'h8079: data_out = 8'h79;
                    16'h807A: data_out = 8'h7A;
                    16'h807B: data_out = 8'h7B;
                    16'h807C: data_out = 8'h7C;
                    16'h807D: data_out = 8'h7D;
                    16'h807E: data_out = 8'h7E;
                    16'h807F: data_out = 8'h7F;
                    16'h8080: data_out = 8'h0;
                    16'h8081: data_out = 8'h81;
                    16'h8082: data_out = 8'h82;
                    16'h8083: data_out = 8'h83;
                    16'h8084: data_out = 8'h84;
                    16'h8085: data_out = 8'h85;
                    16'h8086: data_out = 8'h86;
                    16'h8087: data_out = 8'h87;
                    16'h8088: data_out = 8'h88;
                    16'h8089: data_out = 8'h89;
                    16'h808A: data_out = 8'h8A;
                    16'h808B: data_out = 8'h8B;
                    16'h808C: data_out = 8'h8C;
                    16'h808D: data_out = 8'h8D;
                    16'h808E: data_out = 8'h8E;
                    16'h808F: data_out = 8'h8F;
                    16'h8090: data_out = 8'h90;
                    16'h8091: data_out = 8'h91;
                    16'h8092: data_out = 8'h92;
                    16'h8093: data_out = 8'h93;
                    16'h8094: data_out = 8'h94;
                    16'h8095: data_out = 8'h95;
                    16'h8096: data_out = 8'h96;
                    16'h8097: data_out = 8'h97;
                    16'h8098: data_out = 8'h98;
                    16'h8099: data_out = 8'h99;
                    16'h809A: data_out = 8'h9A;
                    16'h809B: data_out = 8'h9B;
                    16'h809C: data_out = 8'h9C;
                    16'h809D: data_out = 8'h9D;
                    16'h809E: data_out = 8'h9E;
                    16'h809F: data_out = 8'h9F;
                    16'h80A0: data_out = 8'hA0;
                    16'h80A1: data_out = 8'hA1;
                    16'h80A2: data_out = 8'hA2;
                    16'h80A3: data_out = 8'hA3;
                    16'h80A4: data_out = 8'hA4;
                    16'h80A5: data_out = 8'hA5;
                    16'h80A6: data_out = 8'hA6;
                    16'h80A7: data_out = 8'hA7;
                    16'h80A8: data_out = 8'hA8;
                    16'h80A9: data_out = 8'hA9;
                    16'h80AA: data_out = 8'hAA;
                    16'h80AB: data_out = 8'hAB;
                    16'h80AC: data_out = 8'hAC;
                    16'h80AD: data_out = 8'hAD;
                    16'h80AE: data_out = 8'hAE;
                    16'h80AF: data_out = 8'hAF;
                    16'h80B0: data_out = 8'hB0;
                    16'h80B1: data_out = 8'hB1;
                    16'h80B2: data_out = 8'hB2;
                    16'h80B3: data_out = 8'hB3;
                    16'h80B4: data_out = 8'hB4;
                    16'h80B5: data_out = 8'hB5;
                    16'h80B6: data_out = 8'hB6;
                    16'h80B7: data_out = 8'hB7;
                    16'h80B8: data_out = 8'hB8;
                    16'h80B9: data_out = 8'hB9;
                    16'h80BA: data_out = 8'hBA;
                    16'h80BB: data_out = 8'hBB;
                    16'h80BC: data_out = 8'hBC;
                    16'h80BD: data_out = 8'hBD;
                    16'h80BE: data_out = 8'hBE;
                    16'h80BF: data_out = 8'hBF;
                    16'h80C0: data_out = 8'hC0;
                    16'h80C1: data_out = 8'hC1;
                    16'h80C2: data_out = 8'hC2;
                    16'h80C3: data_out = 8'hC3;
                    16'h80C4: data_out = 8'hC4;
                    16'h80C5: data_out = 8'hC5;
                    16'h80C6: data_out = 8'hC6;
                    16'h80C7: data_out = 8'hC7;
                    16'h80C8: data_out = 8'hC8;
                    16'h80C9: data_out = 8'hC9;
                    16'h80CA: data_out = 8'hCA;
                    16'h80CB: data_out = 8'hCB;
                    16'h80CC: data_out = 8'hCC;
                    16'h80CD: data_out = 8'hCD;
                    16'h80CE: data_out = 8'hCE;
                    16'h80CF: data_out = 8'hCF;
                    16'h80D0: data_out = 8'hD0;
                    16'h80D1: data_out = 8'hD1;
                    16'h80D2: data_out = 8'hD2;
                    16'h80D3: data_out = 8'hD3;
                    16'h80D4: data_out = 8'hD4;
                    16'h80D5: data_out = 8'hD5;
                    16'h80D6: data_out = 8'hD6;
                    16'h80D7: data_out = 8'hD7;
                    16'h80D8: data_out = 8'hD8;
                    16'h80D9: data_out = 8'hD9;
                    16'h80DA: data_out = 8'hDA;
                    16'h80DB: data_out = 8'hDB;
                    16'h80DC: data_out = 8'hDC;
                    16'h80DD: data_out = 8'hDD;
                    16'h80DE: data_out = 8'hDE;
                    16'h80DF: data_out = 8'hDF;
                    16'h80E0: data_out = 8'hE0;
                    16'h80E1: data_out = 8'hE1;
                    16'h80E2: data_out = 8'hE2;
                    16'h80E3: data_out = 8'hE3;
                    16'h80E4: data_out = 8'hE4;
                    16'h80E5: data_out = 8'hE5;
                    16'h80E6: data_out = 8'hE6;
                    16'h80E7: data_out = 8'hE7;
                    16'h80E8: data_out = 8'hE8;
                    16'h80E9: data_out = 8'hE9;
                    16'h80EA: data_out = 8'hEA;
                    16'h80EB: data_out = 8'hEB;
                    16'h80EC: data_out = 8'hEC;
                    16'h80ED: data_out = 8'hED;
                    16'h80EE: data_out = 8'hEE;
                    16'h80EF: data_out = 8'hEF;
                    16'h80F0: data_out = 8'hF0;
                    16'h80F1: data_out = 8'hF1;
                    16'h80F2: data_out = 8'hF2;
                    16'h80F3: data_out = 8'hF3;
                    16'h80F4: data_out = 8'hF4;
                    16'h80F5: data_out = 8'hF5;
                    16'h80F6: data_out = 8'hF6;
                    16'h80F7: data_out = 8'hF7;
                    16'h80F8: data_out = 8'hF8;
                    16'h80F9: data_out = 8'hF9;
                    16'h80FA: data_out = 8'hFA;
                    16'h80FB: data_out = 8'hFB;
                    16'h80FC: data_out = 8'hFC;
                    16'h80FD: data_out = 8'hFD;
                    16'h80FE: data_out = 8'hFE;
                    16'h80FF: data_out = 8'hFF;
                    16'h8100: data_out = 8'h81;
                    16'h8101: data_out = 8'h0;
                    16'h8102: data_out = 8'h1;
                    16'h8103: data_out = 8'h2;
                    16'h8104: data_out = 8'h3;
                    16'h8105: data_out = 8'h4;
                    16'h8106: data_out = 8'h5;
                    16'h8107: data_out = 8'h6;
                    16'h8108: data_out = 8'h7;
                    16'h8109: data_out = 8'h8;
                    16'h810A: data_out = 8'h9;
                    16'h810B: data_out = 8'hA;
                    16'h810C: data_out = 8'hB;
                    16'h810D: data_out = 8'hC;
                    16'h810E: data_out = 8'hD;
                    16'h810F: data_out = 8'hE;
                    16'h8110: data_out = 8'hF;
                    16'h8111: data_out = 8'h10;
                    16'h8112: data_out = 8'h11;
                    16'h8113: data_out = 8'h12;
                    16'h8114: data_out = 8'h13;
                    16'h8115: data_out = 8'h14;
                    16'h8116: data_out = 8'h15;
                    16'h8117: data_out = 8'h16;
                    16'h8118: data_out = 8'h17;
                    16'h8119: data_out = 8'h18;
                    16'h811A: data_out = 8'h19;
                    16'h811B: data_out = 8'h1A;
                    16'h811C: data_out = 8'h1B;
                    16'h811D: data_out = 8'h1C;
                    16'h811E: data_out = 8'h1D;
                    16'h811F: data_out = 8'h1E;
                    16'h8120: data_out = 8'h1F;
                    16'h8121: data_out = 8'h20;
                    16'h8122: data_out = 8'h21;
                    16'h8123: data_out = 8'h22;
                    16'h8124: data_out = 8'h23;
                    16'h8125: data_out = 8'h24;
                    16'h8126: data_out = 8'h25;
                    16'h8127: data_out = 8'h26;
                    16'h8128: data_out = 8'h27;
                    16'h8129: data_out = 8'h28;
                    16'h812A: data_out = 8'h29;
                    16'h812B: data_out = 8'h2A;
                    16'h812C: data_out = 8'h2B;
                    16'h812D: data_out = 8'h2C;
                    16'h812E: data_out = 8'h2D;
                    16'h812F: data_out = 8'h2E;
                    16'h8130: data_out = 8'h2F;
                    16'h8131: data_out = 8'h30;
                    16'h8132: data_out = 8'h31;
                    16'h8133: data_out = 8'h32;
                    16'h8134: data_out = 8'h33;
                    16'h8135: data_out = 8'h34;
                    16'h8136: data_out = 8'h35;
                    16'h8137: data_out = 8'h36;
                    16'h8138: data_out = 8'h37;
                    16'h8139: data_out = 8'h38;
                    16'h813A: data_out = 8'h39;
                    16'h813B: data_out = 8'h3A;
                    16'h813C: data_out = 8'h3B;
                    16'h813D: data_out = 8'h3C;
                    16'h813E: data_out = 8'h3D;
                    16'h813F: data_out = 8'h3E;
                    16'h8140: data_out = 8'h3F;
                    16'h8141: data_out = 8'h40;
                    16'h8142: data_out = 8'h41;
                    16'h8143: data_out = 8'h42;
                    16'h8144: data_out = 8'h43;
                    16'h8145: data_out = 8'h44;
                    16'h8146: data_out = 8'h45;
                    16'h8147: data_out = 8'h46;
                    16'h8148: data_out = 8'h47;
                    16'h8149: data_out = 8'h48;
                    16'h814A: data_out = 8'h49;
                    16'h814B: data_out = 8'h4A;
                    16'h814C: data_out = 8'h4B;
                    16'h814D: data_out = 8'h4C;
                    16'h814E: data_out = 8'h4D;
                    16'h814F: data_out = 8'h4E;
                    16'h8150: data_out = 8'h4F;
                    16'h8151: data_out = 8'h50;
                    16'h8152: data_out = 8'h51;
                    16'h8153: data_out = 8'h52;
                    16'h8154: data_out = 8'h53;
                    16'h8155: data_out = 8'h54;
                    16'h8156: data_out = 8'h55;
                    16'h8157: data_out = 8'h56;
                    16'h8158: data_out = 8'h57;
                    16'h8159: data_out = 8'h58;
                    16'h815A: data_out = 8'h59;
                    16'h815B: data_out = 8'h5A;
                    16'h815C: data_out = 8'h5B;
                    16'h815D: data_out = 8'h5C;
                    16'h815E: data_out = 8'h5D;
                    16'h815F: data_out = 8'h5E;
                    16'h8160: data_out = 8'h5F;
                    16'h8161: data_out = 8'h60;
                    16'h8162: data_out = 8'h61;
                    16'h8163: data_out = 8'h62;
                    16'h8164: data_out = 8'h63;
                    16'h8165: data_out = 8'h64;
                    16'h8166: data_out = 8'h65;
                    16'h8167: data_out = 8'h66;
                    16'h8168: data_out = 8'h67;
                    16'h8169: data_out = 8'h68;
                    16'h816A: data_out = 8'h69;
                    16'h816B: data_out = 8'h6A;
                    16'h816C: data_out = 8'h6B;
                    16'h816D: data_out = 8'h6C;
                    16'h816E: data_out = 8'h6D;
                    16'h816F: data_out = 8'h6E;
                    16'h8170: data_out = 8'h6F;
                    16'h8171: data_out = 8'h70;
                    16'h8172: data_out = 8'h71;
                    16'h8173: data_out = 8'h72;
                    16'h8174: data_out = 8'h73;
                    16'h8175: data_out = 8'h74;
                    16'h8176: data_out = 8'h75;
                    16'h8177: data_out = 8'h76;
                    16'h8178: data_out = 8'h77;
                    16'h8179: data_out = 8'h78;
                    16'h817A: data_out = 8'h79;
                    16'h817B: data_out = 8'h7A;
                    16'h817C: data_out = 8'h7B;
                    16'h817D: data_out = 8'h7C;
                    16'h817E: data_out = 8'h7D;
                    16'h817F: data_out = 8'h7E;
                    16'h8180: data_out = 8'h81;
                    16'h8181: data_out = 8'h82;
                    16'h8182: data_out = 8'h83;
                    16'h8183: data_out = 8'h84;
                    16'h8184: data_out = 8'h85;
                    16'h8185: data_out = 8'h86;
                    16'h8186: data_out = 8'h87;
                    16'h8187: data_out = 8'h88;
                    16'h8188: data_out = 8'h89;
                    16'h8189: data_out = 8'h8A;
                    16'h818A: data_out = 8'h8B;
                    16'h818B: data_out = 8'h8C;
                    16'h818C: data_out = 8'h8D;
                    16'h818D: data_out = 8'h8E;
                    16'h818E: data_out = 8'h8F;
                    16'h818F: data_out = 8'h90;
                    16'h8190: data_out = 8'h91;
                    16'h8191: data_out = 8'h92;
                    16'h8192: data_out = 8'h93;
                    16'h8193: data_out = 8'h94;
                    16'h8194: data_out = 8'h95;
                    16'h8195: data_out = 8'h96;
                    16'h8196: data_out = 8'h97;
                    16'h8197: data_out = 8'h98;
                    16'h8198: data_out = 8'h99;
                    16'h8199: data_out = 8'h9A;
                    16'h819A: data_out = 8'h9B;
                    16'h819B: data_out = 8'h9C;
                    16'h819C: data_out = 8'h9D;
                    16'h819D: data_out = 8'h9E;
                    16'h819E: data_out = 8'h9F;
                    16'h819F: data_out = 8'hA0;
                    16'h81A0: data_out = 8'hA1;
                    16'h81A1: data_out = 8'hA2;
                    16'h81A2: data_out = 8'hA3;
                    16'h81A3: data_out = 8'hA4;
                    16'h81A4: data_out = 8'hA5;
                    16'h81A5: data_out = 8'hA6;
                    16'h81A6: data_out = 8'hA7;
                    16'h81A7: data_out = 8'hA8;
                    16'h81A8: data_out = 8'hA9;
                    16'h81A9: data_out = 8'hAA;
                    16'h81AA: data_out = 8'hAB;
                    16'h81AB: data_out = 8'hAC;
                    16'h81AC: data_out = 8'hAD;
                    16'h81AD: data_out = 8'hAE;
                    16'h81AE: data_out = 8'hAF;
                    16'h81AF: data_out = 8'hB0;
                    16'h81B0: data_out = 8'hB1;
                    16'h81B1: data_out = 8'hB2;
                    16'h81B2: data_out = 8'hB3;
                    16'h81B3: data_out = 8'hB4;
                    16'h81B4: data_out = 8'hB5;
                    16'h81B5: data_out = 8'hB6;
                    16'h81B6: data_out = 8'hB7;
                    16'h81B7: data_out = 8'hB8;
                    16'h81B8: data_out = 8'hB9;
                    16'h81B9: data_out = 8'hBA;
                    16'h81BA: data_out = 8'hBB;
                    16'h81BB: data_out = 8'hBC;
                    16'h81BC: data_out = 8'hBD;
                    16'h81BD: data_out = 8'hBE;
                    16'h81BE: data_out = 8'hBF;
                    16'h81BF: data_out = 8'hC0;
                    16'h81C0: data_out = 8'hC1;
                    16'h81C1: data_out = 8'hC2;
                    16'h81C2: data_out = 8'hC3;
                    16'h81C3: data_out = 8'hC4;
                    16'h81C4: data_out = 8'hC5;
                    16'h81C5: data_out = 8'hC6;
                    16'h81C6: data_out = 8'hC7;
                    16'h81C7: data_out = 8'hC8;
                    16'h81C8: data_out = 8'hC9;
                    16'h81C9: data_out = 8'hCA;
                    16'h81CA: data_out = 8'hCB;
                    16'h81CB: data_out = 8'hCC;
                    16'h81CC: data_out = 8'hCD;
                    16'h81CD: data_out = 8'hCE;
                    16'h81CE: data_out = 8'hCF;
                    16'h81CF: data_out = 8'hD0;
                    16'h81D0: data_out = 8'hD1;
                    16'h81D1: data_out = 8'hD2;
                    16'h81D2: data_out = 8'hD3;
                    16'h81D3: data_out = 8'hD4;
                    16'h81D4: data_out = 8'hD5;
                    16'h81D5: data_out = 8'hD6;
                    16'h81D6: data_out = 8'hD7;
                    16'h81D7: data_out = 8'hD8;
                    16'h81D8: data_out = 8'hD9;
                    16'h81D9: data_out = 8'hDA;
                    16'h81DA: data_out = 8'hDB;
                    16'h81DB: data_out = 8'hDC;
                    16'h81DC: data_out = 8'hDD;
                    16'h81DD: data_out = 8'hDE;
                    16'h81DE: data_out = 8'hDF;
                    16'h81DF: data_out = 8'hE0;
                    16'h81E0: data_out = 8'hE1;
                    16'h81E1: data_out = 8'hE2;
                    16'h81E2: data_out = 8'hE3;
                    16'h81E3: data_out = 8'hE4;
                    16'h81E4: data_out = 8'hE5;
                    16'h81E5: data_out = 8'hE6;
                    16'h81E6: data_out = 8'hE7;
                    16'h81E7: data_out = 8'hE8;
                    16'h81E8: data_out = 8'hE9;
                    16'h81E9: data_out = 8'hEA;
                    16'h81EA: data_out = 8'hEB;
                    16'h81EB: data_out = 8'hEC;
                    16'h81EC: data_out = 8'hED;
                    16'h81ED: data_out = 8'hEE;
                    16'h81EE: data_out = 8'hEF;
                    16'h81EF: data_out = 8'hF0;
                    16'h81F0: data_out = 8'hF1;
                    16'h81F1: data_out = 8'hF2;
                    16'h81F2: data_out = 8'hF3;
                    16'h81F3: data_out = 8'hF4;
                    16'h81F4: data_out = 8'hF5;
                    16'h81F5: data_out = 8'hF6;
                    16'h81F6: data_out = 8'hF7;
                    16'h81F7: data_out = 8'hF8;
                    16'h81F8: data_out = 8'hF9;
                    16'h81F9: data_out = 8'hFA;
                    16'h81FA: data_out = 8'hFB;
                    16'h81FB: data_out = 8'hFC;
                    16'h81FC: data_out = 8'hFD;
                    16'h81FD: data_out = 8'hFE;
                    16'h81FE: data_out = 8'hFF;
                    16'h81FF: data_out = 8'h80;
                    16'h8200: data_out = 8'h82;
                    16'h8201: data_out = 8'h81;
                    16'h8202: data_out = 8'h0;
                    16'h8203: data_out = 8'h1;
                    16'h8204: data_out = 8'h2;
                    16'h8205: data_out = 8'h3;
                    16'h8206: data_out = 8'h4;
                    16'h8207: data_out = 8'h5;
                    16'h8208: data_out = 8'h6;
                    16'h8209: data_out = 8'h7;
                    16'h820A: data_out = 8'h8;
                    16'h820B: data_out = 8'h9;
                    16'h820C: data_out = 8'hA;
                    16'h820D: data_out = 8'hB;
                    16'h820E: data_out = 8'hC;
                    16'h820F: data_out = 8'hD;
                    16'h8210: data_out = 8'hE;
                    16'h8211: data_out = 8'hF;
                    16'h8212: data_out = 8'h10;
                    16'h8213: data_out = 8'h11;
                    16'h8214: data_out = 8'h12;
                    16'h8215: data_out = 8'h13;
                    16'h8216: data_out = 8'h14;
                    16'h8217: data_out = 8'h15;
                    16'h8218: data_out = 8'h16;
                    16'h8219: data_out = 8'h17;
                    16'h821A: data_out = 8'h18;
                    16'h821B: data_out = 8'h19;
                    16'h821C: data_out = 8'h1A;
                    16'h821D: data_out = 8'h1B;
                    16'h821E: data_out = 8'h1C;
                    16'h821F: data_out = 8'h1D;
                    16'h8220: data_out = 8'h1E;
                    16'h8221: data_out = 8'h1F;
                    16'h8222: data_out = 8'h20;
                    16'h8223: data_out = 8'h21;
                    16'h8224: data_out = 8'h22;
                    16'h8225: data_out = 8'h23;
                    16'h8226: data_out = 8'h24;
                    16'h8227: data_out = 8'h25;
                    16'h8228: data_out = 8'h26;
                    16'h8229: data_out = 8'h27;
                    16'h822A: data_out = 8'h28;
                    16'h822B: data_out = 8'h29;
                    16'h822C: data_out = 8'h2A;
                    16'h822D: data_out = 8'h2B;
                    16'h822E: data_out = 8'h2C;
                    16'h822F: data_out = 8'h2D;
                    16'h8230: data_out = 8'h2E;
                    16'h8231: data_out = 8'h2F;
                    16'h8232: data_out = 8'h30;
                    16'h8233: data_out = 8'h31;
                    16'h8234: data_out = 8'h32;
                    16'h8235: data_out = 8'h33;
                    16'h8236: data_out = 8'h34;
                    16'h8237: data_out = 8'h35;
                    16'h8238: data_out = 8'h36;
                    16'h8239: data_out = 8'h37;
                    16'h823A: data_out = 8'h38;
                    16'h823B: data_out = 8'h39;
                    16'h823C: data_out = 8'h3A;
                    16'h823D: data_out = 8'h3B;
                    16'h823E: data_out = 8'h3C;
                    16'h823F: data_out = 8'h3D;
                    16'h8240: data_out = 8'h3E;
                    16'h8241: data_out = 8'h3F;
                    16'h8242: data_out = 8'h40;
                    16'h8243: data_out = 8'h41;
                    16'h8244: data_out = 8'h42;
                    16'h8245: data_out = 8'h43;
                    16'h8246: data_out = 8'h44;
                    16'h8247: data_out = 8'h45;
                    16'h8248: data_out = 8'h46;
                    16'h8249: data_out = 8'h47;
                    16'h824A: data_out = 8'h48;
                    16'h824B: data_out = 8'h49;
                    16'h824C: data_out = 8'h4A;
                    16'h824D: data_out = 8'h4B;
                    16'h824E: data_out = 8'h4C;
                    16'h824F: data_out = 8'h4D;
                    16'h8250: data_out = 8'h4E;
                    16'h8251: data_out = 8'h4F;
                    16'h8252: data_out = 8'h50;
                    16'h8253: data_out = 8'h51;
                    16'h8254: data_out = 8'h52;
                    16'h8255: data_out = 8'h53;
                    16'h8256: data_out = 8'h54;
                    16'h8257: data_out = 8'h55;
                    16'h8258: data_out = 8'h56;
                    16'h8259: data_out = 8'h57;
                    16'h825A: data_out = 8'h58;
                    16'h825B: data_out = 8'h59;
                    16'h825C: data_out = 8'h5A;
                    16'h825D: data_out = 8'h5B;
                    16'h825E: data_out = 8'h5C;
                    16'h825F: data_out = 8'h5D;
                    16'h8260: data_out = 8'h5E;
                    16'h8261: data_out = 8'h5F;
                    16'h8262: data_out = 8'h60;
                    16'h8263: data_out = 8'h61;
                    16'h8264: data_out = 8'h62;
                    16'h8265: data_out = 8'h63;
                    16'h8266: data_out = 8'h64;
                    16'h8267: data_out = 8'h65;
                    16'h8268: data_out = 8'h66;
                    16'h8269: data_out = 8'h67;
                    16'h826A: data_out = 8'h68;
                    16'h826B: data_out = 8'h69;
                    16'h826C: data_out = 8'h6A;
                    16'h826D: data_out = 8'h6B;
                    16'h826E: data_out = 8'h6C;
                    16'h826F: data_out = 8'h6D;
                    16'h8270: data_out = 8'h6E;
                    16'h8271: data_out = 8'h6F;
                    16'h8272: data_out = 8'h70;
                    16'h8273: data_out = 8'h71;
                    16'h8274: data_out = 8'h72;
                    16'h8275: data_out = 8'h73;
                    16'h8276: data_out = 8'h74;
                    16'h8277: data_out = 8'h75;
                    16'h8278: data_out = 8'h76;
                    16'h8279: data_out = 8'h77;
                    16'h827A: data_out = 8'h78;
                    16'h827B: data_out = 8'h79;
                    16'h827C: data_out = 8'h7A;
                    16'h827D: data_out = 8'h7B;
                    16'h827E: data_out = 8'h7C;
                    16'h827F: data_out = 8'h7D;
                    16'h8280: data_out = 8'h82;
                    16'h8281: data_out = 8'h83;
                    16'h8282: data_out = 8'h84;
                    16'h8283: data_out = 8'h85;
                    16'h8284: data_out = 8'h86;
                    16'h8285: data_out = 8'h87;
                    16'h8286: data_out = 8'h88;
                    16'h8287: data_out = 8'h89;
                    16'h8288: data_out = 8'h8A;
                    16'h8289: data_out = 8'h8B;
                    16'h828A: data_out = 8'h8C;
                    16'h828B: data_out = 8'h8D;
                    16'h828C: data_out = 8'h8E;
                    16'h828D: data_out = 8'h8F;
                    16'h828E: data_out = 8'h90;
                    16'h828F: data_out = 8'h91;
                    16'h8290: data_out = 8'h92;
                    16'h8291: data_out = 8'h93;
                    16'h8292: data_out = 8'h94;
                    16'h8293: data_out = 8'h95;
                    16'h8294: data_out = 8'h96;
                    16'h8295: data_out = 8'h97;
                    16'h8296: data_out = 8'h98;
                    16'h8297: data_out = 8'h99;
                    16'h8298: data_out = 8'h9A;
                    16'h8299: data_out = 8'h9B;
                    16'h829A: data_out = 8'h9C;
                    16'h829B: data_out = 8'h9D;
                    16'h829C: data_out = 8'h9E;
                    16'h829D: data_out = 8'h9F;
                    16'h829E: data_out = 8'hA0;
                    16'h829F: data_out = 8'hA1;
                    16'h82A0: data_out = 8'hA2;
                    16'h82A1: data_out = 8'hA3;
                    16'h82A2: data_out = 8'hA4;
                    16'h82A3: data_out = 8'hA5;
                    16'h82A4: data_out = 8'hA6;
                    16'h82A5: data_out = 8'hA7;
                    16'h82A6: data_out = 8'hA8;
                    16'h82A7: data_out = 8'hA9;
                    16'h82A8: data_out = 8'hAA;
                    16'h82A9: data_out = 8'hAB;
                    16'h82AA: data_out = 8'hAC;
                    16'h82AB: data_out = 8'hAD;
                    16'h82AC: data_out = 8'hAE;
                    16'h82AD: data_out = 8'hAF;
                    16'h82AE: data_out = 8'hB0;
                    16'h82AF: data_out = 8'hB1;
                    16'h82B0: data_out = 8'hB2;
                    16'h82B1: data_out = 8'hB3;
                    16'h82B2: data_out = 8'hB4;
                    16'h82B3: data_out = 8'hB5;
                    16'h82B4: data_out = 8'hB6;
                    16'h82B5: data_out = 8'hB7;
                    16'h82B6: data_out = 8'hB8;
                    16'h82B7: data_out = 8'hB9;
                    16'h82B8: data_out = 8'hBA;
                    16'h82B9: data_out = 8'hBB;
                    16'h82BA: data_out = 8'hBC;
                    16'h82BB: data_out = 8'hBD;
                    16'h82BC: data_out = 8'hBE;
                    16'h82BD: data_out = 8'hBF;
                    16'h82BE: data_out = 8'hC0;
                    16'h82BF: data_out = 8'hC1;
                    16'h82C0: data_out = 8'hC2;
                    16'h82C1: data_out = 8'hC3;
                    16'h82C2: data_out = 8'hC4;
                    16'h82C3: data_out = 8'hC5;
                    16'h82C4: data_out = 8'hC6;
                    16'h82C5: data_out = 8'hC7;
                    16'h82C6: data_out = 8'hC8;
                    16'h82C7: data_out = 8'hC9;
                    16'h82C8: data_out = 8'hCA;
                    16'h82C9: data_out = 8'hCB;
                    16'h82CA: data_out = 8'hCC;
                    16'h82CB: data_out = 8'hCD;
                    16'h82CC: data_out = 8'hCE;
                    16'h82CD: data_out = 8'hCF;
                    16'h82CE: data_out = 8'hD0;
                    16'h82CF: data_out = 8'hD1;
                    16'h82D0: data_out = 8'hD2;
                    16'h82D1: data_out = 8'hD3;
                    16'h82D2: data_out = 8'hD4;
                    16'h82D3: data_out = 8'hD5;
                    16'h82D4: data_out = 8'hD6;
                    16'h82D5: data_out = 8'hD7;
                    16'h82D6: data_out = 8'hD8;
                    16'h82D7: data_out = 8'hD9;
                    16'h82D8: data_out = 8'hDA;
                    16'h82D9: data_out = 8'hDB;
                    16'h82DA: data_out = 8'hDC;
                    16'h82DB: data_out = 8'hDD;
                    16'h82DC: data_out = 8'hDE;
                    16'h82DD: data_out = 8'hDF;
                    16'h82DE: data_out = 8'hE0;
                    16'h82DF: data_out = 8'hE1;
                    16'h82E0: data_out = 8'hE2;
                    16'h82E1: data_out = 8'hE3;
                    16'h82E2: data_out = 8'hE4;
                    16'h82E3: data_out = 8'hE5;
                    16'h82E4: data_out = 8'hE6;
                    16'h82E5: data_out = 8'hE7;
                    16'h82E6: data_out = 8'hE8;
                    16'h82E7: data_out = 8'hE9;
                    16'h82E8: data_out = 8'hEA;
                    16'h82E9: data_out = 8'hEB;
                    16'h82EA: data_out = 8'hEC;
                    16'h82EB: data_out = 8'hED;
                    16'h82EC: data_out = 8'hEE;
                    16'h82ED: data_out = 8'hEF;
                    16'h82EE: data_out = 8'hF0;
                    16'h82EF: data_out = 8'hF1;
                    16'h82F0: data_out = 8'hF2;
                    16'h82F1: data_out = 8'hF3;
                    16'h82F2: data_out = 8'hF4;
                    16'h82F3: data_out = 8'hF5;
                    16'h82F4: data_out = 8'hF6;
                    16'h82F5: data_out = 8'hF7;
                    16'h82F6: data_out = 8'hF8;
                    16'h82F7: data_out = 8'hF9;
                    16'h82F8: data_out = 8'hFA;
                    16'h82F9: data_out = 8'hFB;
                    16'h82FA: data_out = 8'hFC;
                    16'h82FB: data_out = 8'hFD;
                    16'h82FC: data_out = 8'hFE;
                    16'h82FD: data_out = 8'hFF;
                    16'h82FE: data_out = 8'h80;
                    16'h82FF: data_out = 8'h81;
                    16'h8300: data_out = 8'h83;
                    16'h8301: data_out = 8'h82;
                    16'h8302: data_out = 8'h81;
                    16'h8303: data_out = 8'h0;
                    16'h8304: data_out = 8'h1;
                    16'h8305: data_out = 8'h2;
                    16'h8306: data_out = 8'h3;
                    16'h8307: data_out = 8'h4;
                    16'h8308: data_out = 8'h5;
                    16'h8309: data_out = 8'h6;
                    16'h830A: data_out = 8'h7;
                    16'h830B: data_out = 8'h8;
                    16'h830C: data_out = 8'h9;
                    16'h830D: data_out = 8'hA;
                    16'h830E: data_out = 8'hB;
                    16'h830F: data_out = 8'hC;
                    16'h8310: data_out = 8'hD;
                    16'h8311: data_out = 8'hE;
                    16'h8312: data_out = 8'hF;
                    16'h8313: data_out = 8'h10;
                    16'h8314: data_out = 8'h11;
                    16'h8315: data_out = 8'h12;
                    16'h8316: data_out = 8'h13;
                    16'h8317: data_out = 8'h14;
                    16'h8318: data_out = 8'h15;
                    16'h8319: data_out = 8'h16;
                    16'h831A: data_out = 8'h17;
                    16'h831B: data_out = 8'h18;
                    16'h831C: data_out = 8'h19;
                    16'h831D: data_out = 8'h1A;
                    16'h831E: data_out = 8'h1B;
                    16'h831F: data_out = 8'h1C;
                    16'h8320: data_out = 8'h1D;
                    16'h8321: data_out = 8'h1E;
                    16'h8322: data_out = 8'h1F;
                    16'h8323: data_out = 8'h20;
                    16'h8324: data_out = 8'h21;
                    16'h8325: data_out = 8'h22;
                    16'h8326: data_out = 8'h23;
                    16'h8327: data_out = 8'h24;
                    16'h8328: data_out = 8'h25;
                    16'h8329: data_out = 8'h26;
                    16'h832A: data_out = 8'h27;
                    16'h832B: data_out = 8'h28;
                    16'h832C: data_out = 8'h29;
                    16'h832D: data_out = 8'h2A;
                    16'h832E: data_out = 8'h2B;
                    16'h832F: data_out = 8'h2C;
                    16'h8330: data_out = 8'h2D;
                    16'h8331: data_out = 8'h2E;
                    16'h8332: data_out = 8'h2F;
                    16'h8333: data_out = 8'h30;
                    16'h8334: data_out = 8'h31;
                    16'h8335: data_out = 8'h32;
                    16'h8336: data_out = 8'h33;
                    16'h8337: data_out = 8'h34;
                    16'h8338: data_out = 8'h35;
                    16'h8339: data_out = 8'h36;
                    16'h833A: data_out = 8'h37;
                    16'h833B: data_out = 8'h38;
                    16'h833C: data_out = 8'h39;
                    16'h833D: data_out = 8'h3A;
                    16'h833E: data_out = 8'h3B;
                    16'h833F: data_out = 8'h3C;
                    16'h8340: data_out = 8'h3D;
                    16'h8341: data_out = 8'h3E;
                    16'h8342: data_out = 8'h3F;
                    16'h8343: data_out = 8'h40;
                    16'h8344: data_out = 8'h41;
                    16'h8345: data_out = 8'h42;
                    16'h8346: data_out = 8'h43;
                    16'h8347: data_out = 8'h44;
                    16'h8348: data_out = 8'h45;
                    16'h8349: data_out = 8'h46;
                    16'h834A: data_out = 8'h47;
                    16'h834B: data_out = 8'h48;
                    16'h834C: data_out = 8'h49;
                    16'h834D: data_out = 8'h4A;
                    16'h834E: data_out = 8'h4B;
                    16'h834F: data_out = 8'h4C;
                    16'h8350: data_out = 8'h4D;
                    16'h8351: data_out = 8'h4E;
                    16'h8352: data_out = 8'h4F;
                    16'h8353: data_out = 8'h50;
                    16'h8354: data_out = 8'h51;
                    16'h8355: data_out = 8'h52;
                    16'h8356: data_out = 8'h53;
                    16'h8357: data_out = 8'h54;
                    16'h8358: data_out = 8'h55;
                    16'h8359: data_out = 8'h56;
                    16'h835A: data_out = 8'h57;
                    16'h835B: data_out = 8'h58;
                    16'h835C: data_out = 8'h59;
                    16'h835D: data_out = 8'h5A;
                    16'h835E: data_out = 8'h5B;
                    16'h835F: data_out = 8'h5C;
                    16'h8360: data_out = 8'h5D;
                    16'h8361: data_out = 8'h5E;
                    16'h8362: data_out = 8'h5F;
                    16'h8363: data_out = 8'h60;
                    16'h8364: data_out = 8'h61;
                    16'h8365: data_out = 8'h62;
                    16'h8366: data_out = 8'h63;
                    16'h8367: data_out = 8'h64;
                    16'h8368: data_out = 8'h65;
                    16'h8369: data_out = 8'h66;
                    16'h836A: data_out = 8'h67;
                    16'h836B: data_out = 8'h68;
                    16'h836C: data_out = 8'h69;
                    16'h836D: data_out = 8'h6A;
                    16'h836E: data_out = 8'h6B;
                    16'h836F: data_out = 8'h6C;
                    16'h8370: data_out = 8'h6D;
                    16'h8371: data_out = 8'h6E;
                    16'h8372: data_out = 8'h6F;
                    16'h8373: data_out = 8'h70;
                    16'h8374: data_out = 8'h71;
                    16'h8375: data_out = 8'h72;
                    16'h8376: data_out = 8'h73;
                    16'h8377: data_out = 8'h74;
                    16'h8378: data_out = 8'h75;
                    16'h8379: data_out = 8'h76;
                    16'h837A: data_out = 8'h77;
                    16'h837B: data_out = 8'h78;
                    16'h837C: data_out = 8'h79;
                    16'h837D: data_out = 8'h7A;
                    16'h837E: data_out = 8'h7B;
                    16'h837F: data_out = 8'h7C;
                    16'h8380: data_out = 8'h83;
                    16'h8381: data_out = 8'h84;
                    16'h8382: data_out = 8'h85;
                    16'h8383: data_out = 8'h86;
                    16'h8384: data_out = 8'h87;
                    16'h8385: data_out = 8'h88;
                    16'h8386: data_out = 8'h89;
                    16'h8387: data_out = 8'h8A;
                    16'h8388: data_out = 8'h8B;
                    16'h8389: data_out = 8'h8C;
                    16'h838A: data_out = 8'h8D;
                    16'h838B: data_out = 8'h8E;
                    16'h838C: data_out = 8'h8F;
                    16'h838D: data_out = 8'h90;
                    16'h838E: data_out = 8'h91;
                    16'h838F: data_out = 8'h92;
                    16'h8390: data_out = 8'h93;
                    16'h8391: data_out = 8'h94;
                    16'h8392: data_out = 8'h95;
                    16'h8393: data_out = 8'h96;
                    16'h8394: data_out = 8'h97;
                    16'h8395: data_out = 8'h98;
                    16'h8396: data_out = 8'h99;
                    16'h8397: data_out = 8'h9A;
                    16'h8398: data_out = 8'h9B;
                    16'h8399: data_out = 8'h9C;
                    16'h839A: data_out = 8'h9D;
                    16'h839B: data_out = 8'h9E;
                    16'h839C: data_out = 8'h9F;
                    16'h839D: data_out = 8'hA0;
                    16'h839E: data_out = 8'hA1;
                    16'h839F: data_out = 8'hA2;
                    16'h83A0: data_out = 8'hA3;
                    16'h83A1: data_out = 8'hA4;
                    16'h83A2: data_out = 8'hA5;
                    16'h83A3: data_out = 8'hA6;
                    16'h83A4: data_out = 8'hA7;
                    16'h83A5: data_out = 8'hA8;
                    16'h83A6: data_out = 8'hA9;
                    16'h83A7: data_out = 8'hAA;
                    16'h83A8: data_out = 8'hAB;
                    16'h83A9: data_out = 8'hAC;
                    16'h83AA: data_out = 8'hAD;
                    16'h83AB: data_out = 8'hAE;
                    16'h83AC: data_out = 8'hAF;
                    16'h83AD: data_out = 8'hB0;
                    16'h83AE: data_out = 8'hB1;
                    16'h83AF: data_out = 8'hB2;
                    16'h83B0: data_out = 8'hB3;
                    16'h83B1: data_out = 8'hB4;
                    16'h83B2: data_out = 8'hB5;
                    16'h83B3: data_out = 8'hB6;
                    16'h83B4: data_out = 8'hB7;
                    16'h83B5: data_out = 8'hB8;
                    16'h83B6: data_out = 8'hB9;
                    16'h83B7: data_out = 8'hBA;
                    16'h83B8: data_out = 8'hBB;
                    16'h83B9: data_out = 8'hBC;
                    16'h83BA: data_out = 8'hBD;
                    16'h83BB: data_out = 8'hBE;
                    16'h83BC: data_out = 8'hBF;
                    16'h83BD: data_out = 8'hC0;
                    16'h83BE: data_out = 8'hC1;
                    16'h83BF: data_out = 8'hC2;
                    16'h83C0: data_out = 8'hC3;
                    16'h83C1: data_out = 8'hC4;
                    16'h83C2: data_out = 8'hC5;
                    16'h83C3: data_out = 8'hC6;
                    16'h83C4: data_out = 8'hC7;
                    16'h83C5: data_out = 8'hC8;
                    16'h83C6: data_out = 8'hC9;
                    16'h83C7: data_out = 8'hCA;
                    16'h83C8: data_out = 8'hCB;
                    16'h83C9: data_out = 8'hCC;
                    16'h83CA: data_out = 8'hCD;
                    16'h83CB: data_out = 8'hCE;
                    16'h83CC: data_out = 8'hCF;
                    16'h83CD: data_out = 8'hD0;
                    16'h83CE: data_out = 8'hD1;
                    16'h83CF: data_out = 8'hD2;
                    16'h83D0: data_out = 8'hD3;
                    16'h83D1: data_out = 8'hD4;
                    16'h83D2: data_out = 8'hD5;
                    16'h83D3: data_out = 8'hD6;
                    16'h83D4: data_out = 8'hD7;
                    16'h83D5: data_out = 8'hD8;
                    16'h83D6: data_out = 8'hD9;
                    16'h83D7: data_out = 8'hDA;
                    16'h83D8: data_out = 8'hDB;
                    16'h83D9: data_out = 8'hDC;
                    16'h83DA: data_out = 8'hDD;
                    16'h83DB: data_out = 8'hDE;
                    16'h83DC: data_out = 8'hDF;
                    16'h83DD: data_out = 8'hE0;
                    16'h83DE: data_out = 8'hE1;
                    16'h83DF: data_out = 8'hE2;
                    16'h83E0: data_out = 8'hE3;
                    16'h83E1: data_out = 8'hE4;
                    16'h83E2: data_out = 8'hE5;
                    16'h83E3: data_out = 8'hE6;
                    16'h83E4: data_out = 8'hE7;
                    16'h83E5: data_out = 8'hE8;
                    16'h83E6: data_out = 8'hE9;
                    16'h83E7: data_out = 8'hEA;
                    16'h83E8: data_out = 8'hEB;
                    16'h83E9: data_out = 8'hEC;
                    16'h83EA: data_out = 8'hED;
                    16'h83EB: data_out = 8'hEE;
                    16'h83EC: data_out = 8'hEF;
                    16'h83ED: data_out = 8'hF0;
                    16'h83EE: data_out = 8'hF1;
                    16'h83EF: data_out = 8'hF2;
                    16'h83F0: data_out = 8'hF3;
                    16'h83F1: data_out = 8'hF4;
                    16'h83F2: data_out = 8'hF5;
                    16'h83F3: data_out = 8'hF6;
                    16'h83F4: data_out = 8'hF7;
                    16'h83F5: data_out = 8'hF8;
                    16'h83F6: data_out = 8'hF9;
                    16'h83F7: data_out = 8'hFA;
                    16'h83F8: data_out = 8'hFB;
                    16'h83F9: data_out = 8'hFC;
                    16'h83FA: data_out = 8'hFD;
                    16'h83FB: data_out = 8'hFE;
                    16'h83FC: data_out = 8'hFF;
                    16'h83FD: data_out = 8'h80;
                    16'h83FE: data_out = 8'h81;
                    16'h83FF: data_out = 8'h82;
                    16'h8400: data_out = 8'h84;
                    16'h8401: data_out = 8'h83;
                    16'h8402: data_out = 8'h82;
                    16'h8403: data_out = 8'h81;
                    16'h8404: data_out = 8'h0;
                    16'h8405: data_out = 8'h1;
                    16'h8406: data_out = 8'h2;
                    16'h8407: data_out = 8'h3;
                    16'h8408: data_out = 8'h4;
                    16'h8409: data_out = 8'h5;
                    16'h840A: data_out = 8'h6;
                    16'h840B: data_out = 8'h7;
                    16'h840C: data_out = 8'h8;
                    16'h840D: data_out = 8'h9;
                    16'h840E: data_out = 8'hA;
                    16'h840F: data_out = 8'hB;
                    16'h8410: data_out = 8'hC;
                    16'h8411: data_out = 8'hD;
                    16'h8412: data_out = 8'hE;
                    16'h8413: data_out = 8'hF;
                    16'h8414: data_out = 8'h10;
                    16'h8415: data_out = 8'h11;
                    16'h8416: data_out = 8'h12;
                    16'h8417: data_out = 8'h13;
                    16'h8418: data_out = 8'h14;
                    16'h8419: data_out = 8'h15;
                    16'h841A: data_out = 8'h16;
                    16'h841B: data_out = 8'h17;
                    16'h841C: data_out = 8'h18;
                    16'h841D: data_out = 8'h19;
                    16'h841E: data_out = 8'h1A;
                    16'h841F: data_out = 8'h1B;
                    16'h8420: data_out = 8'h1C;
                    16'h8421: data_out = 8'h1D;
                    16'h8422: data_out = 8'h1E;
                    16'h8423: data_out = 8'h1F;
                    16'h8424: data_out = 8'h20;
                    16'h8425: data_out = 8'h21;
                    16'h8426: data_out = 8'h22;
                    16'h8427: data_out = 8'h23;
                    16'h8428: data_out = 8'h24;
                    16'h8429: data_out = 8'h25;
                    16'h842A: data_out = 8'h26;
                    16'h842B: data_out = 8'h27;
                    16'h842C: data_out = 8'h28;
                    16'h842D: data_out = 8'h29;
                    16'h842E: data_out = 8'h2A;
                    16'h842F: data_out = 8'h2B;
                    16'h8430: data_out = 8'h2C;
                    16'h8431: data_out = 8'h2D;
                    16'h8432: data_out = 8'h2E;
                    16'h8433: data_out = 8'h2F;
                    16'h8434: data_out = 8'h30;
                    16'h8435: data_out = 8'h31;
                    16'h8436: data_out = 8'h32;
                    16'h8437: data_out = 8'h33;
                    16'h8438: data_out = 8'h34;
                    16'h8439: data_out = 8'h35;
                    16'h843A: data_out = 8'h36;
                    16'h843B: data_out = 8'h37;
                    16'h843C: data_out = 8'h38;
                    16'h843D: data_out = 8'h39;
                    16'h843E: data_out = 8'h3A;
                    16'h843F: data_out = 8'h3B;
                    16'h8440: data_out = 8'h3C;
                    16'h8441: data_out = 8'h3D;
                    16'h8442: data_out = 8'h3E;
                    16'h8443: data_out = 8'h3F;
                    16'h8444: data_out = 8'h40;
                    16'h8445: data_out = 8'h41;
                    16'h8446: data_out = 8'h42;
                    16'h8447: data_out = 8'h43;
                    16'h8448: data_out = 8'h44;
                    16'h8449: data_out = 8'h45;
                    16'h844A: data_out = 8'h46;
                    16'h844B: data_out = 8'h47;
                    16'h844C: data_out = 8'h48;
                    16'h844D: data_out = 8'h49;
                    16'h844E: data_out = 8'h4A;
                    16'h844F: data_out = 8'h4B;
                    16'h8450: data_out = 8'h4C;
                    16'h8451: data_out = 8'h4D;
                    16'h8452: data_out = 8'h4E;
                    16'h8453: data_out = 8'h4F;
                    16'h8454: data_out = 8'h50;
                    16'h8455: data_out = 8'h51;
                    16'h8456: data_out = 8'h52;
                    16'h8457: data_out = 8'h53;
                    16'h8458: data_out = 8'h54;
                    16'h8459: data_out = 8'h55;
                    16'h845A: data_out = 8'h56;
                    16'h845B: data_out = 8'h57;
                    16'h845C: data_out = 8'h58;
                    16'h845D: data_out = 8'h59;
                    16'h845E: data_out = 8'h5A;
                    16'h845F: data_out = 8'h5B;
                    16'h8460: data_out = 8'h5C;
                    16'h8461: data_out = 8'h5D;
                    16'h8462: data_out = 8'h5E;
                    16'h8463: data_out = 8'h5F;
                    16'h8464: data_out = 8'h60;
                    16'h8465: data_out = 8'h61;
                    16'h8466: data_out = 8'h62;
                    16'h8467: data_out = 8'h63;
                    16'h8468: data_out = 8'h64;
                    16'h8469: data_out = 8'h65;
                    16'h846A: data_out = 8'h66;
                    16'h846B: data_out = 8'h67;
                    16'h846C: data_out = 8'h68;
                    16'h846D: data_out = 8'h69;
                    16'h846E: data_out = 8'h6A;
                    16'h846F: data_out = 8'h6B;
                    16'h8470: data_out = 8'h6C;
                    16'h8471: data_out = 8'h6D;
                    16'h8472: data_out = 8'h6E;
                    16'h8473: data_out = 8'h6F;
                    16'h8474: data_out = 8'h70;
                    16'h8475: data_out = 8'h71;
                    16'h8476: data_out = 8'h72;
                    16'h8477: data_out = 8'h73;
                    16'h8478: data_out = 8'h74;
                    16'h8479: data_out = 8'h75;
                    16'h847A: data_out = 8'h76;
                    16'h847B: data_out = 8'h77;
                    16'h847C: data_out = 8'h78;
                    16'h847D: data_out = 8'h79;
                    16'h847E: data_out = 8'h7A;
                    16'h847F: data_out = 8'h7B;
                    16'h8480: data_out = 8'h84;
                    16'h8481: data_out = 8'h85;
                    16'h8482: data_out = 8'h86;
                    16'h8483: data_out = 8'h87;
                    16'h8484: data_out = 8'h88;
                    16'h8485: data_out = 8'h89;
                    16'h8486: data_out = 8'h8A;
                    16'h8487: data_out = 8'h8B;
                    16'h8488: data_out = 8'h8C;
                    16'h8489: data_out = 8'h8D;
                    16'h848A: data_out = 8'h8E;
                    16'h848B: data_out = 8'h8F;
                    16'h848C: data_out = 8'h90;
                    16'h848D: data_out = 8'h91;
                    16'h848E: data_out = 8'h92;
                    16'h848F: data_out = 8'h93;
                    16'h8490: data_out = 8'h94;
                    16'h8491: data_out = 8'h95;
                    16'h8492: data_out = 8'h96;
                    16'h8493: data_out = 8'h97;
                    16'h8494: data_out = 8'h98;
                    16'h8495: data_out = 8'h99;
                    16'h8496: data_out = 8'h9A;
                    16'h8497: data_out = 8'h9B;
                    16'h8498: data_out = 8'h9C;
                    16'h8499: data_out = 8'h9D;
                    16'h849A: data_out = 8'h9E;
                    16'h849B: data_out = 8'h9F;
                    16'h849C: data_out = 8'hA0;
                    16'h849D: data_out = 8'hA1;
                    16'h849E: data_out = 8'hA2;
                    16'h849F: data_out = 8'hA3;
                    16'h84A0: data_out = 8'hA4;
                    16'h84A1: data_out = 8'hA5;
                    16'h84A2: data_out = 8'hA6;
                    16'h84A3: data_out = 8'hA7;
                    16'h84A4: data_out = 8'hA8;
                    16'h84A5: data_out = 8'hA9;
                    16'h84A6: data_out = 8'hAA;
                    16'h84A7: data_out = 8'hAB;
                    16'h84A8: data_out = 8'hAC;
                    16'h84A9: data_out = 8'hAD;
                    16'h84AA: data_out = 8'hAE;
                    16'h84AB: data_out = 8'hAF;
                    16'h84AC: data_out = 8'hB0;
                    16'h84AD: data_out = 8'hB1;
                    16'h84AE: data_out = 8'hB2;
                    16'h84AF: data_out = 8'hB3;
                    16'h84B0: data_out = 8'hB4;
                    16'h84B1: data_out = 8'hB5;
                    16'h84B2: data_out = 8'hB6;
                    16'h84B3: data_out = 8'hB7;
                    16'h84B4: data_out = 8'hB8;
                    16'h84B5: data_out = 8'hB9;
                    16'h84B6: data_out = 8'hBA;
                    16'h84B7: data_out = 8'hBB;
                    16'h84B8: data_out = 8'hBC;
                    16'h84B9: data_out = 8'hBD;
                    16'h84BA: data_out = 8'hBE;
                    16'h84BB: data_out = 8'hBF;
                    16'h84BC: data_out = 8'hC0;
                    16'h84BD: data_out = 8'hC1;
                    16'h84BE: data_out = 8'hC2;
                    16'h84BF: data_out = 8'hC3;
                    16'h84C0: data_out = 8'hC4;
                    16'h84C1: data_out = 8'hC5;
                    16'h84C2: data_out = 8'hC6;
                    16'h84C3: data_out = 8'hC7;
                    16'h84C4: data_out = 8'hC8;
                    16'h84C5: data_out = 8'hC9;
                    16'h84C6: data_out = 8'hCA;
                    16'h84C7: data_out = 8'hCB;
                    16'h84C8: data_out = 8'hCC;
                    16'h84C9: data_out = 8'hCD;
                    16'h84CA: data_out = 8'hCE;
                    16'h84CB: data_out = 8'hCF;
                    16'h84CC: data_out = 8'hD0;
                    16'h84CD: data_out = 8'hD1;
                    16'h84CE: data_out = 8'hD2;
                    16'h84CF: data_out = 8'hD3;
                    16'h84D0: data_out = 8'hD4;
                    16'h84D1: data_out = 8'hD5;
                    16'h84D2: data_out = 8'hD6;
                    16'h84D3: data_out = 8'hD7;
                    16'h84D4: data_out = 8'hD8;
                    16'h84D5: data_out = 8'hD9;
                    16'h84D6: data_out = 8'hDA;
                    16'h84D7: data_out = 8'hDB;
                    16'h84D8: data_out = 8'hDC;
                    16'h84D9: data_out = 8'hDD;
                    16'h84DA: data_out = 8'hDE;
                    16'h84DB: data_out = 8'hDF;
                    16'h84DC: data_out = 8'hE0;
                    16'h84DD: data_out = 8'hE1;
                    16'h84DE: data_out = 8'hE2;
                    16'h84DF: data_out = 8'hE3;
                    16'h84E0: data_out = 8'hE4;
                    16'h84E1: data_out = 8'hE5;
                    16'h84E2: data_out = 8'hE6;
                    16'h84E3: data_out = 8'hE7;
                    16'h84E4: data_out = 8'hE8;
                    16'h84E5: data_out = 8'hE9;
                    16'h84E6: data_out = 8'hEA;
                    16'h84E7: data_out = 8'hEB;
                    16'h84E8: data_out = 8'hEC;
                    16'h84E9: data_out = 8'hED;
                    16'h84EA: data_out = 8'hEE;
                    16'h84EB: data_out = 8'hEF;
                    16'h84EC: data_out = 8'hF0;
                    16'h84ED: data_out = 8'hF1;
                    16'h84EE: data_out = 8'hF2;
                    16'h84EF: data_out = 8'hF3;
                    16'h84F0: data_out = 8'hF4;
                    16'h84F1: data_out = 8'hF5;
                    16'h84F2: data_out = 8'hF6;
                    16'h84F3: data_out = 8'hF7;
                    16'h84F4: data_out = 8'hF8;
                    16'h84F5: data_out = 8'hF9;
                    16'h84F6: data_out = 8'hFA;
                    16'h84F7: data_out = 8'hFB;
                    16'h84F8: data_out = 8'hFC;
                    16'h84F9: data_out = 8'hFD;
                    16'h84FA: data_out = 8'hFE;
                    16'h84FB: data_out = 8'hFF;
                    16'h84FC: data_out = 8'h80;
                    16'h84FD: data_out = 8'h81;
                    16'h84FE: data_out = 8'h82;
                    16'h84FF: data_out = 8'h83;
                    16'h8500: data_out = 8'h85;
                    16'h8501: data_out = 8'h84;
                    16'h8502: data_out = 8'h83;
                    16'h8503: data_out = 8'h82;
                    16'h8504: data_out = 8'h81;
                    16'h8505: data_out = 8'h0;
                    16'h8506: data_out = 8'h1;
                    16'h8507: data_out = 8'h2;
                    16'h8508: data_out = 8'h3;
                    16'h8509: data_out = 8'h4;
                    16'h850A: data_out = 8'h5;
                    16'h850B: data_out = 8'h6;
                    16'h850C: data_out = 8'h7;
                    16'h850D: data_out = 8'h8;
                    16'h850E: data_out = 8'h9;
                    16'h850F: data_out = 8'hA;
                    16'h8510: data_out = 8'hB;
                    16'h8511: data_out = 8'hC;
                    16'h8512: data_out = 8'hD;
                    16'h8513: data_out = 8'hE;
                    16'h8514: data_out = 8'hF;
                    16'h8515: data_out = 8'h10;
                    16'h8516: data_out = 8'h11;
                    16'h8517: data_out = 8'h12;
                    16'h8518: data_out = 8'h13;
                    16'h8519: data_out = 8'h14;
                    16'h851A: data_out = 8'h15;
                    16'h851B: data_out = 8'h16;
                    16'h851C: data_out = 8'h17;
                    16'h851D: data_out = 8'h18;
                    16'h851E: data_out = 8'h19;
                    16'h851F: data_out = 8'h1A;
                    16'h8520: data_out = 8'h1B;
                    16'h8521: data_out = 8'h1C;
                    16'h8522: data_out = 8'h1D;
                    16'h8523: data_out = 8'h1E;
                    16'h8524: data_out = 8'h1F;
                    16'h8525: data_out = 8'h20;
                    16'h8526: data_out = 8'h21;
                    16'h8527: data_out = 8'h22;
                    16'h8528: data_out = 8'h23;
                    16'h8529: data_out = 8'h24;
                    16'h852A: data_out = 8'h25;
                    16'h852B: data_out = 8'h26;
                    16'h852C: data_out = 8'h27;
                    16'h852D: data_out = 8'h28;
                    16'h852E: data_out = 8'h29;
                    16'h852F: data_out = 8'h2A;
                    16'h8530: data_out = 8'h2B;
                    16'h8531: data_out = 8'h2C;
                    16'h8532: data_out = 8'h2D;
                    16'h8533: data_out = 8'h2E;
                    16'h8534: data_out = 8'h2F;
                    16'h8535: data_out = 8'h30;
                    16'h8536: data_out = 8'h31;
                    16'h8537: data_out = 8'h32;
                    16'h8538: data_out = 8'h33;
                    16'h8539: data_out = 8'h34;
                    16'h853A: data_out = 8'h35;
                    16'h853B: data_out = 8'h36;
                    16'h853C: data_out = 8'h37;
                    16'h853D: data_out = 8'h38;
                    16'h853E: data_out = 8'h39;
                    16'h853F: data_out = 8'h3A;
                    16'h8540: data_out = 8'h3B;
                    16'h8541: data_out = 8'h3C;
                    16'h8542: data_out = 8'h3D;
                    16'h8543: data_out = 8'h3E;
                    16'h8544: data_out = 8'h3F;
                    16'h8545: data_out = 8'h40;
                    16'h8546: data_out = 8'h41;
                    16'h8547: data_out = 8'h42;
                    16'h8548: data_out = 8'h43;
                    16'h8549: data_out = 8'h44;
                    16'h854A: data_out = 8'h45;
                    16'h854B: data_out = 8'h46;
                    16'h854C: data_out = 8'h47;
                    16'h854D: data_out = 8'h48;
                    16'h854E: data_out = 8'h49;
                    16'h854F: data_out = 8'h4A;
                    16'h8550: data_out = 8'h4B;
                    16'h8551: data_out = 8'h4C;
                    16'h8552: data_out = 8'h4D;
                    16'h8553: data_out = 8'h4E;
                    16'h8554: data_out = 8'h4F;
                    16'h8555: data_out = 8'h50;
                    16'h8556: data_out = 8'h51;
                    16'h8557: data_out = 8'h52;
                    16'h8558: data_out = 8'h53;
                    16'h8559: data_out = 8'h54;
                    16'h855A: data_out = 8'h55;
                    16'h855B: data_out = 8'h56;
                    16'h855C: data_out = 8'h57;
                    16'h855D: data_out = 8'h58;
                    16'h855E: data_out = 8'h59;
                    16'h855F: data_out = 8'h5A;
                    16'h8560: data_out = 8'h5B;
                    16'h8561: data_out = 8'h5C;
                    16'h8562: data_out = 8'h5D;
                    16'h8563: data_out = 8'h5E;
                    16'h8564: data_out = 8'h5F;
                    16'h8565: data_out = 8'h60;
                    16'h8566: data_out = 8'h61;
                    16'h8567: data_out = 8'h62;
                    16'h8568: data_out = 8'h63;
                    16'h8569: data_out = 8'h64;
                    16'h856A: data_out = 8'h65;
                    16'h856B: data_out = 8'h66;
                    16'h856C: data_out = 8'h67;
                    16'h856D: data_out = 8'h68;
                    16'h856E: data_out = 8'h69;
                    16'h856F: data_out = 8'h6A;
                    16'h8570: data_out = 8'h6B;
                    16'h8571: data_out = 8'h6C;
                    16'h8572: data_out = 8'h6D;
                    16'h8573: data_out = 8'h6E;
                    16'h8574: data_out = 8'h6F;
                    16'h8575: data_out = 8'h70;
                    16'h8576: data_out = 8'h71;
                    16'h8577: data_out = 8'h72;
                    16'h8578: data_out = 8'h73;
                    16'h8579: data_out = 8'h74;
                    16'h857A: data_out = 8'h75;
                    16'h857B: data_out = 8'h76;
                    16'h857C: data_out = 8'h77;
                    16'h857D: data_out = 8'h78;
                    16'h857E: data_out = 8'h79;
                    16'h857F: data_out = 8'h7A;
                    16'h8580: data_out = 8'h85;
                    16'h8581: data_out = 8'h86;
                    16'h8582: data_out = 8'h87;
                    16'h8583: data_out = 8'h88;
                    16'h8584: data_out = 8'h89;
                    16'h8585: data_out = 8'h8A;
                    16'h8586: data_out = 8'h8B;
                    16'h8587: data_out = 8'h8C;
                    16'h8588: data_out = 8'h8D;
                    16'h8589: data_out = 8'h8E;
                    16'h858A: data_out = 8'h8F;
                    16'h858B: data_out = 8'h90;
                    16'h858C: data_out = 8'h91;
                    16'h858D: data_out = 8'h92;
                    16'h858E: data_out = 8'h93;
                    16'h858F: data_out = 8'h94;
                    16'h8590: data_out = 8'h95;
                    16'h8591: data_out = 8'h96;
                    16'h8592: data_out = 8'h97;
                    16'h8593: data_out = 8'h98;
                    16'h8594: data_out = 8'h99;
                    16'h8595: data_out = 8'h9A;
                    16'h8596: data_out = 8'h9B;
                    16'h8597: data_out = 8'h9C;
                    16'h8598: data_out = 8'h9D;
                    16'h8599: data_out = 8'h9E;
                    16'h859A: data_out = 8'h9F;
                    16'h859B: data_out = 8'hA0;
                    16'h859C: data_out = 8'hA1;
                    16'h859D: data_out = 8'hA2;
                    16'h859E: data_out = 8'hA3;
                    16'h859F: data_out = 8'hA4;
                    16'h85A0: data_out = 8'hA5;
                    16'h85A1: data_out = 8'hA6;
                    16'h85A2: data_out = 8'hA7;
                    16'h85A3: data_out = 8'hA8;
                    16'h85A4: data_out = 8'hA9;
                    16'h85A5: data_out = 8'hAA;
                    16'h85A6: data_out = 8'hAB;
                    16'h85A7: data_out = 8'hAC;
                    16'h85A8: data_out = 8'hAD;
                    16'h85A9: data_out = 8'hAE;
                    16'h85AA: data_out = 8'hAF;
                    16'h85AB: data_out = 8'hB0;
                    16'h85AC: data_out = 8'hB1;
                    16'h85AD: data_out = 8'hB2;
                    16'h85AE: data_out = 8'hB3;
                    16'h85AF: data_out = 8'hB4;
                    16'h85B0: data_out = 8'hB5;
                    16'h85B1: data_out = 8'hB6;
                    16'h85B2: data_out = 8'hB7;
                    16'h85B3: data_out = 8'hB8;
                    16'h85B4: data_out = 8'hB9;
                    16'h85B5: data_out = 8'hBA;
                    16'h85B6: data_out = 8'hBB;
                    16'h85B7: data_out = 8'hBC;
                    16'h85B8: data_out = 8'hBD;
                    16'h85B9: data_out = 8'hBE;
                    16'h85BA: data_out = 8'hBF;
                    16'h85BB: data_out = 8'hC0;
                    16'h85BC: data_out = 8'hC1;
                    16'h85BD: data_out = 8'hC2;
                    16'h85BE: data_out = 8'hC3;
                    16'h85BF: data_out = 8'hC4;
                    16'h85C0: data_out = 8'hC5;
                    16'h85C1: data_out = 8'hC6;
                    16'h85C2: data_out = 8'hC7;
                    16'h85C3: data_out = 8'hC8;
                    16'h85C4: data_out = 8'hC9;
                    16'h85C5: data_out = 8'hCA;
                    16'h85C6: data_out = 8'hCB;
                    16'h85C7: data_out = 8'hCC;
                    16'h85C8: data_out = 8'hCD;
                    16'h85C9: data_out = 8'hCE;
                    16'h85CA: data_out = 8'hCF;
                    16'h85CB: data_out = 8'hD0;
                    16'h85CC: data_out = 8'hD1;
                    16'h85CD: data_out = 8'hD2;
                    16'h85CE: data_out = 8'hD3;
                    16'h85CF: data_out = 8'hD4;
                    16'h85D0: data_out = 8'hD5;
                    16'h85D1: data_out = 8'hD6;
                    16'h85D2: data_out = 8'hD7;
                    16'h85D3: data_out = 8'hD8;
                    16'h85D4: data_out = 8'hD9;
                    16'h85D5: data_out = 8'hDA;
                    16'h85D6: data_out = 8'hDB;
                    16'h85D7: data_out = 8'hDC;
                    16'h85D8: data_out = 8'hDD;
                    16'h85D9: data_out = 8'hDE;
                    16'h85DA: data_out = 8'hDF;
                    16'h85DB: data_out = 8'hE0;
                    16'h85DC: data_out = 8'hE1;
                    16'h85DD: data_out = 8'hE2;
                    16'h85DE: data_out = 8'hE3;
                    16'h85DF: data_out = 8'hE4;
                    16'h85E0: data_out = 8'hE5;
                    16'h85E1: data_out = 8'hE6;
                    16'h85E2: data_out = 8'hE7;
                    16'h85E3: data_out = 8'hE8;
                    16'h85E4: data_out = 8'hE9;
                    16'h85E5: data_out = 8'hEA;
                    16'h85E6: data_out = 8'hEB;
                    16'h85E7: data_out = 8'hEC;
                    16'h85E8: data_out = 8'hED;
                    16'h85E9: data_out = 8'hEE;
                    16'h85EA: data_out = 8'hEF;
                    16'h85EB: data_out = 8'hF0;
                    16'h85EC: data_out = 8'hF1;
                    16'h85ED: data_out = 8'hF2;
                    16'h85EE: data_out = 8'hF3;
                    16'h85EF: data_out = 8'hF4;
                    16'h85F0: data_out = 8'hF5;
                    16'h85F1: data_out = 8'hF6;
                    16'h85F2: data_out = 8'hF7;
                    16'h85F3: data_out = 8'hF8;
                    16'h85F4: data_out = 8'hF9;
                    16'h85F5: data_out = 8'hFA;
                    16'h85F6: data_out = 8'hFB;
                    16'h85F7: data_out = 8'hFC;
                    16'h85F8: data_out = 8'hFD;
                    16'h85F9: data_out = 8'hFE;
                    16'h85FA: data_out = 8'hFF;
                    16'h85FB: data_out = 8'h80;
                    16'h85FC: data_out = 8'h81;
                    16'h85FD: data_out = 8'h82;
                    16'h85FE: data_out = 8'h83;
                    16'h85FF: data_out = 8'h84;
                    16'h8600: data_out = 8'h86;
                    16'h8601: data_out = 8'h85;
                    16'h8602: data_out = 8'h84;
                    16'h8603: data_out = 8'h83;
                    16'h8604: data_out = 8'h82;
                    16'h8605: data_out = 8'h81;
                    16'h8606: data_out = 8'h0;
                    16'h8607: data_out = 8'h1;
                    16'h8608: data_out = 8'h2;
                    16'h8609: data_out = 8'h3;
                    16'h860A: data_out = 8'h4;
                    16'h860B: data_out = 8'h5;
                    16'h860C: data_out = 8'h6;
                    16'h860D: data_out = 8'h7;
                    16'h860E: data_out = 8'h8;
                    16'h860F: data_out = 8'h9;
                    16'h8610: data_out = 8'hA;
                    16'h8611: data_out = 8'hB;
                    16'h8612: data_out = 8'hC;
                    16'h8613: data_out = 8'hD;
                    16'h8614: data_out = 8'hE;
                    16'h8615: data_out = 8'hF;
                    16'h8616: data_out = 8'h10;
                    16'h8617: data_out = 8'h11;
                    16'h8618: data_out = 8'h12;
                    16'h8619: data_out = 8'h13;
                    16'h861A: data_out = 8'h14;
                    16'h861B: data_out = 8'h15;
                    16'h861C: data_out = 8'h16;
                    16'h861D: data_out = 8'h17;
                    16'h861E: data_out = 8'h18;
                    16'h861F: data_out = 8'h19;
                    16'h8620: data_out = 8'h1A;
                    16'h8621: data_out = 8'h1B;
                    16'h8622: data_out = 8'h1C;
                    16'h8623: data_out = 8'h1D;
                    16'h8624: data_out = 8'h1E;
                    16'h8625: data_out = 8'h1F;
                    16'h8626: data_out = 8'h20;
                    16'h8627: data_out = 8'h21;
                    16'h8628: data_out = 8'h22;
                    16'h8629: data_out = 8'h23;
                    16'h862A: data_out = 8'h24;
                    16'h862B: data_out = 8'h25;
                    16'h862C: data_out = 8'h26;
                    16'h862D: data_out = 8'h27;
                    16'h862E: data_out = 8'h28;
                    16'h862F: data_out = 8'h29;
                    16'h8630: data_out = 8'h2A;
                    16'h8631: data_out = 8'h2B;
                    16'h8632: data_out = 8'h2C;
                    16'h8633: data_out = 8'h2D;
                    16'h8634: data_out = 8'h2E;
                    16'h8635: data_out = 8'h2F;
                    16'h8636: data_out = 8'h30;
                    16'h8637: data_out = 8'h31;
                    16'h8638: data_out = 8'h32;
                    16'h8639: data_out = 8'h33;
                    16'h863A: data_out = 8'h34;
                    16'h863B: data_out = 8'h35;
                    16'h863C: data_out = 8'h36;
                    16'h863D: data_out = 8'h37;
                    16'h863E: data_out = 8'h38;
                    16'h863F: data_out = 8'h39;
                    16'h8640: data_out = 8'h3A;
                    16'h8641: data_out = 8'h3B;
                    16'h8642: data_out = 8'h3C;
                    16'h8643: data_out = 8'h3D;
                    16'h8644: data_out = 8'h3E;
                    16'h8645: data_out = 8'h3F;
                    16'h8646: data_out = 8'h40;
                    16'h8647: data_out = 8'h41;
                    16'h8648: data_out = 8'h42;
                    16'h8649: data_out = 8'h43;
                    16'h864A: data_out = 8'h44;
                    16'h864B: data_out = 8'h45;
                    16'h864C: data_out = 8'h46;
                    16'h864D: data_out = 8'h47;
                    16'h864E: data_out = 8'h48;
                    16'h864F: data_out = 8'h49;
                    16'h8650: data_out = 8'h4A;
                    16'h8651: data_out = 8'h4B;
                    16'h8652: data_out = 8'h4C;
                    16'h8653: data_out = 8'h4D;
                    16'h8654: data_out = 8'h4E;
                    16'h8655: data_out = 8'h4F;
                    16'h8656: data_out = 8'h50;
                    16'h8657: data_out = 8'h51;
                    16'h8658: data_out = 8'h52;
                    16'h8659: data_out = 8'h53;
                    16'h865A: data_out = 8'h54;
                    16'h865B: data_out = 8'h55;
                    16'h865C: data_out = 8'h56;
                    16'h865D: data_out = 8'h57;
                    16'h865E: data_out = 8'h58;
                    16'h865F: data_out = 8'h59;
                    16'h8660: data_out = 8'h5A;
                    16'h8661: data_out = 8'h5B;
                    16'h8662: data_out = 8'h5C;
                    16'h8663: data_out = 8'h5D;
                    16'h8664: data_out = 8'h5E;
                    16'h8665: data_out = 8'h5F;
                    16'h8666: data_out = 8'h60;
                    16'h8667: data_out = 8'h61;
                    16'h8668: data_out = 8'h62;
                    16'h8669: data_out = 8'h63;
                    16'h866A: data_out = 8'h64;
                    16'h866B: data_out = 8'h65;
                    16'h866C: data_out = 8'h66;
                    16'h866D: data_out = 8'h67;
                    16'h866E: data_out = 8'h68;
                    16'h866F: data_out = 8'h69;
                    16'h8670: data_out = 8'h6A;
                    16'h8671: data_out = 8'h6B;
                    16'h8672: data_out = 8'h6C;
                    16'h8673: data_out = 8'h6D;
                    16'h8674: data_out = 8'h6E;
                    16'h8675: data_out = 8'h6F;
                    16'h8676: data_out = 8'h70;
                    16'h8677: data_out = 8'h71;
                    16'h8678: data_out = 8'h72;
                    16'h8679: data_out = 8'h73;
                    16'h867A: data_out = 8'h74;
                    16'h867B: data_out = 8'h75;
                    16'h867C: data_out = 8'h76;
                    16'h867D: data_out = 8'h77;
                    16'h867E: data_out = 8'h78;
                    16'h867F: data_out = 8'h79;
                    16'h8680: data_out = 8'h86;
                    16'h8681: data_out = 8'h87;
                    16'h8682: data_out = 8'h88;
                    16'h8683: data_out = 8'h89;
                    16'h8684: data_out = 8'h8A;
                    16'h8685: data_out = 8'h8B;
                    16'h8686: data_out = 8'h8C;
                    16'h8687: data_out = 8'h8D;
                    16'h8688: data_out = 8'h8E;
                    16'h8689: data_out = 8'h8F;
                    16'h868A: data_out = 8'h90;
                    16'h868B: data_out = 8'h91;
                    16'h868C: data_out = 8'h92;
                    16'h868D: data_out = 8'h93;
                    16'h868E: data_out = 8'h94;
                    16'h868F: data_out = 8'h95;
                    16'h8690: data_out = 8'h96;
                    16'h8691: data_out = 8'h97;
                    16'h8692: data_out = 8'h98;
                    16'h8693: data_out = 8'h99;
                    16'h8694: data_out = 8'h9A;
                    16'h8695: data_out = 8'h9B;
                    16'h8696: data_out = 8'h9C;
                    16'h8697: data_out = 8'h9D;
                    16'h8698: data_out = 8'h9E;
                    16'h8699: data_out = 8'h9F;
                    16'h869A: data_out = 8'hA0;
                    16'h869B: data_out = 8'hA1;
                    16'h869C: data_out = 8'hA2;
                    16'h869D: data_out = 8'hA3;
                    16'h869E: data_out = 8'hA4;
                    16'h869F: data_out = 8'hA5;
                    16'h86A0: data_out = 8'hA6;
                    16'h86A1: data_out = 8'hA7;
                    16'h86A2: data_out = 8'hA8;
                    16'h86A3: data_out = 8'hA9;
                    16'h86A4: data_out = 8'hAA;
                    16'h86A5: data_out = 8'hAB;
                    16'h86A6: data_out = 8'hAC;
                    16'h86A7: data_out = 8'hAD;
                    16'h86A8: data_out = 8'hAE;
                    16'h86A9: data_out = 8'hAF;
                    16'h86AA: data_out = 8'hB0;
                    16'h86AB: data_out = 8'hB1;
                    16'h86AC: data_out = 8'hB2;
                    16'h86AD: data_out = 8'hB3;
                    16'h86AE: data_out = 8'hB4;
                    16'h86AF: data_out = 8'hB5;
                    16'h86B0: data_out = 8'hB6;
                    16'h86B1: data_out = 8'hB7;
                    16'h86B2: data_out = 8'hB8;
                    16'h86B3: data_out = 8'hB9;
                    16'h86B4: data_out = 8'hBA;
                    16'h86B5: data_out = 8'hBB;
                    16'h86B6: data_out = 8'hBC;
                    16'h86B7: data_out = 8'hBD;
                    16'h86B8: data_out = 8'hBE;
                    16'h86B9: data_out = 8'hBF;
                    16'h86BA: data_out = 8'hC0;
                    16'h86BB: data_out = 8'hC1;
                    16'h86BC: data_out = 8'hC2;
                    16'h86BD: data_out = 8'hC3;
                    16'h86BE: data_out = 8'hC4;
                    16'h86BF: data_out = 8'hC5;
                    16'h86C0: data_out = 8'hC6;
                    16'h86C1: data_out = 8'hC7;
                    16'h86C2: data_out = 8'hC8;
                    16'h86C3: data_out = 8'hC9;
                    16'h86C4: data_out = 8'hCA;
                    16'h86C5: data_out = 8'hCB;
                    16'h86C6: data_out = 8'hCC;
                    16'h86C7: data_out = 8'hCD;
                    16'h86C8: data_out = 8'hCE;
                    16'h86C9: data_out = 8'hCF;
                    16'h86CA: data_out = 8'hD0;
                    16'h86CB: data_out = 8'hD1;
                    16'h86CC: data_out = 8'hD2;
                    16'h86CD: data_out = 8'hD3;
                    16'h86CE: data_out = 8'hD4;
                    16'h86CF: data_out = 8'hD5;
                    16'h86D0: data_out = 8'hD6;
                    16'h86D1: data_out = 8'hD7;
                    16'h86D2: data_out = 8'hD8;
                    16'h86D3: data_out = 8'hD9;
                    16'h86D4: data_out = 8'hDA;
                    16'h86D5: data_out = 8'hDB;
                    16'h86D6: data_out = 8'hDC;
                    16'h86D7: data_out = 8'hDD;
                    16'h86D8: data_out = 8'hDE;
                    16'h86D9: data_out = 8'hDF;
                    16'h86DA: data_out = 8'hE0;
                    16'h86DB: data_out = 8'hE1;
                    16'h86DC: data_out = 8'hE2;
                    16'h86DD: data_out = 8'hE3;
                    16'h86DE: data_out = 8'hE4;
                    16'h86DF: data_out = 8'hE5;
                    16'h86E0: data_out = 8'hE6;
                    16'h86E1: data_out = 8'hE7;
                    16'h86E2: data_out = 8'hE8;
                    16'h86E3: data_out = 8'hE9;
                    16'h86E4: data_out = 8'hEA;
                    16'h86E5: data_out = 8'hEB;
                    16'h86E6: data_out = 8'hEC;
                    16'h86E7: data_out = 8'hED;
                    16'h86E8: data_out = 8'hEE;
                    16'h86E9: data_out = 8'hEF;
                    16'h86EA: data_out = 8'hF0;
                    16'h86EB: data_out = 8'hF1;
                    16'h86EC: data_out = 8'hF2;
                    16'h86ED: data_out = 8'hF3;
                    16'h86EE: data_out = 8'hF4;
                    16'h86EF: data_out = 8'hF5;
                    16'h86F0: data_out = 8'hF6;
                    16'h86F1: data_out = 8'hF7;
                    16'h86F2: data_out = 8'hF8;
                    16'h86F3: data_out = 8'hF9;
                    16'h86F4: data_out = 8'hFA;
                    16'h86F5: data_out = 8'hFB;
                    16'h86F6: data_out = 8'hFC;
                    16'h86F7: data_out = 8'hFD;
                    16'h86F8: data_out = 8'hFE;
                    16'h86F9: data_out = 8'hFF;
                    16'h86FA: data_out = 8'h80;
                    16'h86FB: data_out = 8'h81;
                    16'h86FC: data_out = 8'h82;
                    16'h86FD: data_out = 8'h83;
                    16'h86FE: data_out = 8'h84;
                    16'h86FF: data_out = 8'h85;
                    16'h8700: data_out = 8'h87;
                    16'h8701: data_out = 8'h86;
                    16'h8702: data_out = 8'h85;
                    16'h8703: data_out = 8'h84;
                    16'h8704: data_out = 8'h83;
                    16'h8705: data_out = 8'h82;
                    16'h8706: data_out = 8'h81;
                    16'h8707: data_out = 8'h0;
                    16'h8708: data_out = 8'h1;
                    16'h8709: data_out = 8'h2;
                    16'h870A: data_out = 8'h3;
                    16'h870B: data_out = 8'h4;
                    16'h870C: data_out = 8'h5;
                    16'h870D: data_out = 8'h6;
                    16'h870E: data_out = 8'h7;
                    16'h870F: data_out = 8'h8;
                    16'h8710: data_out = 8'h9;
                    16'h8711: data_out = 8'hA;
                    16'h8712: data_out = 8'hB;
                    16'h8713: data_out = 8'hC;
                    16'h8714: data_out = 8'hD;
                    16'h8715: data_out = 8'hE;
                    16'h8716: data_out = 8'hF;
                    16'h8717: data_out = 8'h10;
                    16'h8718: data_out = 8'h11;
                    16'h8719: data_out = 8'h12;
                    16'h871A: data_out = 8'h13;
                    16'h871B: data_out = 8'h14;
                    16'h871C: data_out = 8'h15;
                    16'h871D: data_out = 8'h16;
                    16'h871E: data_out = 8'h17;
                    16'h871F: data_out = 8'h18;
                    16'h8720: data_out = 8'h19;
                    16'h8721: data_out = 8'h1A;
                    16'h8722: data_out = 8'h1B;
                    16'h8723: data_out = 8'h1C;
                    16'h8724: data_out = 8'h1D;
                    16'h8725: data_out = 8'h1E;
                    16'h8726: data_out = 8'h1F;
                    16'h8727: data_out = 8'h20;
                    16'h8728: data_out = 8'h21;
                    16'h8729: data_out = 8'h22;
                    16'h872A: data_out = 8'h23;
                    16'h872B: data_out = 8'h24;
                    16'h872C: data_out = 8'h25;
                    16'h872D: data_out = 8'h26;
                    16'h872E: data_out = 8'h27;
                    16'h872F: data_out = 8'h28;
                    16'h8730: data_out = 8'h29;
                    16'h8731: data_out = 8'h2A;
                    16'h8732: data_out = 8'h2B;
                    16'h8733: data_out = 8'h2C;
                    16'h8734: data_out = 8'h2D;
                    16'h8735: data_out = 8'h2E;
                    16'h8736: data_out = 8'h2F;
                    16'h8737: data_out = 8'h30;
                    16'h8738: data_out = 8'h31;
                    16'h8739: data_out = 8'h32;
                    16'h873A: data_out = 8'h33;
                    16'h873B: data_out = 8'h34;
                    16'h873C: data_out = 8'h35;
                    16'h873D: data_out = 8'h36;
                    16'h873E: data_out = 8'h37;
                    16'h873F: data_out = 8'h38;
                    16'h8740: data_out = 8'h39;
                    16'h8741: data_out = 8'h3A;
                    16'h8742: data_out = 8'h3B;
                    16'h8743: data_out = 8'h3C;
                    16'h8744: data_out = 8'h3D;
                    16'h8745: data_out = 8'h3E;
                    16'h8746: data_out = 8'h3F;
                    16'h8747: data_out = 8'h40;
                    16'h8748: data_out = 8'h41;
                    16'h8749: data_out = 8'h42;
                    16'h874A: data_out = 8'h43;
                    16'h874B: data_out = 8'h44;
                    16'h874C: data_out = 8'h45;
                    16'h874D: data_out = 8'h46;
                    16'h874E: data_out = 8'h47;
                    16'h874F: data_out = 8'h48;
                    16'h8750: data_out = 8'h49;
                    16'h8751: data_out = 8'h4A;
                    16'h8752: data_out = 8'h4B;
                    16'h8753: data_out = 8'h4C;
                    16'h8754: data_out = 8'h4D;
                    16'h8755: data_out = 8'h4E;
                    16'h8756: data_out = 8'h4F;
                    16'h8757: data_out = 8'h50;
                    16'h8758: data_out = 8'h51;
                    16'h8759: data_out = 8'h52;
                    16'h875A: data_out = 8'h53;
                    16'h875B: data_out = 8'h54;
                    16'h875C: data_out = 8'h55;
                    16'h875D: data_out = 8'h56;
                    16'h875E: data_out = 8'h57;
                    16'h875F: data_out = 8'h58;
                    16'h8760: data_out = 8'h59;
                    16'h8761: data_out = 8'h5A;
                    16'h8762: data_out = 8'h5B;
                    16'h8763: data_out = 8'h5C;
                    16'h8764: data_out = 8'h5D;
                    16'h8765: data_out = 8'h5E;
                    16'h8766: data_out = 8'h5F;
                    16'h8767: data_out = 8'h60;
                    16'h8768: data_out = 8'h61;
                    16'h8769: data_out = 8'h62;
                    16'h876A: data_out = 8'h63;
                    16'h876B: data_out = 8'h64;
                    16'h876C: data_out = 8'h65;
                    16'h876D: data_out = 8'h66;
                    16'h876E: data_out = 8'h67;
                    16'h876F: data_out = 8'h68;
                    16'h8770: data_out = 8'h69;
                    16'h8771: data_out = 8'h6A;
                    16'h8772: data_out = 8'h6B;
                    16'h8773: data_out = 8'h6C;
                    16'h8774: data_out = 8'h6D;
                    16'h8775: data_out = 8'h6E;
                    16'h8776: data_out = 8'h6F;
                    16'h8777: data_out = 8'h70;
                    16'h8778: data_out = 8'h71;
                    16'h8779: data_out = 8'h72;
                    16'h877A: data_out = 8'h73;
                    16'h877B: data_out = 8'h74;
                    16'h877C: data_out = 8'h75;
                    16'h877D: data_out = 8'h76;
                    16'h877E: data_out = 8'h77;
                    16'h877F: data_out = 8'h78;
                    16'h8780: data_out = 8'h87;
                    16'h8781: data_out = 8'h88;
                    16'h8782: data_out = 8'h89;
                    16'h8783: data_out = 8'h8A;
                    16'h8784: data_out = 8'h8B;
                    16'h8785: data_out = 8'h8C;
                    16'h8786: data_out = 8'h8D;
                    16'h8787: data_out = 8'h8E;
                    16'h8788: data_out = 8'h8F;
                    16'h8789: data_out = 8'h90;
                    16'h878A: data_out = 8'h91;
                    16'h878B: data_out = 8'h92;
                    16'h878C: data_out = 8'h93;
                    16'h878D: data_out = 8'h94;
                    16'h878E: data_out = 8'h95;
                    16'h878F: data_out = 8'h96;
                    16'h8790: data_out = 8'h97;
                    16'h8791: data_out = 8'h98;
                    16'h8792: data_out = 8'h99;
                    16'h8793: data_out = 8'h9A;
                    16'h8794: data_out = 8'h9B;
                    16'h8795: data_out = 8'h9C;
                    16'h8796: data_out = 8'h9D;
                    16'h8797: data_out = 8'h9E;
                    16'h8798: data_out = 8'h9F;
                    16'h8799: data_out = 8'hA0;
                    16'h879A: data_out = 8'hA1;
                    16'h879B: data_out = 8'hA2;
                    16'h879C: data_out = 8'hA3;
                    16'h879D: data_out = 8'hA4;
                    16'h879E: data_out = 8'hA5;
                    16'h879F: data_out = 8'hA6;
                    16'h87A0: data_out = 8'hA7;
                    16'h87A1: data_out = 8'hA8;
                    16'h87A2: data_out = 8'hA9;
                    16'h87A3: data_out = 8'hAA;
                    16'h87A4: data_out = 8'hAB;
                    16'h87A5: data_out = 8'hAC;
                    16'h87A6: data_out = 8'hAD;
                    16'h87A7: data_out = 8'hAE;
                    16'h87A8: data_out = 8'hAF;
                    16'h87A9: data_out = 8'hB0;
                    16'h87AA: data_out = 8'hB1;
                    16'h87AB: data_out = 8'hB2;
                    16'h87AC: data_out = 8'hB3;
                    16'h87AD: data_out = 8'hB4;
                    16'h87AE: data_out = 8'hB5;
                    16'h87AF: data_out = 8'hB6;
                    16'h87B0: data_out = 8'hB7;
                    16'h87B1: data_out = 8'hB8;
                    16'h87B2: data_out = 8'hB9;
                    16'h87B3: data_out = 8'hBA;
                    16'h87B4: data_out = 8'hBB;
                    16'h87B5: data_out = 8'hBC;
                    16'h87B6: data_out = 8'hBD;
                    16'h87B7: data_out = 8'hBE;
                    16'h87B8: data_out = 8'hBF;
                    16'h87B9: data_out = 8'hC0;
                    16'h87BA: data_out = 8'hC1;
                    16'h87BB: data_out = 8'hC2;
                    16'h87BC: data_out = 8'hC3;
                    16'h87BD: data_out = 8'hC4;
                    16'h87BE: data_out = 8'hC5;
                    16'h87BF: data_out = 8'hC6;
                    16'h87C0: data_out = 8'hC7;
                    16'h87C1: data_out = 8'hC8;
                    16'h87C2: data_out = 8'hC9;
                    16'h87C3: data_out = 8'hCA;
                    16'h87C4: data_out = 8'hCB;
                    16'h87C5: data_out = 8'hCC;
                    16'h87C6: data_out = 8'hCD;
                    16'h87C7: data_out = 8'hCE;
                    16'h87C8: data_out = 8'hCF;
                    16'h87C9: data_out = 8'hD0;
                    16'h87CA: data_out = 8'hD1;
                    16'h87CB: data_out = 8'hD2;
                    16'h87CC: data_out = 8'hD3;
                    16'h87CD: data_out = 8'hD4;
                    16'h87CE: data_out = 8'hD5;
                    16'h87CF: data_out = 8'hD6;
                    16'h87D0: data_out = 8'hD7;
                    16'h87D1: data_out = 8'hD8;
                    16'h87D2: data_out = 8'hD9;
                    16'h87D3: data_out = 8'hDA;
                    16'h87D4: data_out = 8'hDB;
                    16'h87D5: data_out = 8'hDC;
                    16'h87D6: data_out = 8'hDD;
                    16'h87D7: data_out = 8'hDE;
                    16'h87D8: data_out = 8'hDF;
                    16'h87D9: data_out = 8'hE0;
                    16'h87DA: data_out = 8'hE1;
                    16'h87DB: data_out = 8'hE2;
                    16'h87DC: data_out = 8'hE3;
                    16'h87DD: data_out = 8'hE4;
                    16'h87DE: data_out = 8'hE5;
                    16'h87DF: data_out = 8'hE6;
                    16'h87E0: data_out = 8'hE7;
                    16'h87E1: data_out = 8'hE8;
                    16'h87E2: data_out = 8'hE9;
                    16'h87E3: data_out = 8'hEA;
                    16'h87E4: data_out = 8'hEB;
                    16'h87E5: data_out = 8'hEC;
                    16'h87E6: data_out = 8'hED;
                    16'h87E7: data_out = 8'hEE;
                    16'h87E8: data_out = 8'hEF;
                    16'h87E9: data_out = 8'hF0;
                    16'h87EA: data_out = 8'hF1;
                    16'h87EB: data_out = 8'hF2;
                    16'h87EC: data_out = 8'hF3;
                    16'h87ED: data_out = 8'hF4;
                    16'h87EE: data_out = 8'hF5;
                    16'h87EF: data_out = 8'hF6;
                    16'h87F0: data_out = 8'hF7;
                    16'h87F1: data_out = 8'hF8;
                    16'h87F2: data_out = 8'hF9;
                    16'h87F3: data_out = 8'hFA;
                    16'h87F4: data_out = 8'hFB;
                    16'h87F5: data_out = 8'hFC;
                    16'h87F6: data_out = 8'hFD;
                    16'h87F7: data_out = 8'hFE;
                    16'h87F8: data_out = 8'hFF;
                    16'h87F9: data_out = 8'h80;
                    16'h87FA: data_out = 8'h81;
                    16'h87FB: data_out = 8'h82;
                    16'h87FC: data_out = 8'h83;
                    16'h87FD: data_out = 8'h84;
                    16'h87FE: data_out = 8'h85;
                    16'h87FF: data_out = 8'h86;
                    16'h8800: data_out = 8'h88;
                    16'h8801: data_out = 8'h87;
                    16'h8802: data_out = 8'h86;
                    16'h8803: data_out = 8'h85;
                    16'h8804: data_out = 8'h84;
                    16'h8805: data_out = 8'h83;
                    16'h8806: data_out = 8'h82;
                    16'h8807: data_out = 8'h81;
                    16'h8808: data_out = 8'h0;
                    16'h8809: data_out = 8'h1;
                    16'h880A: data_out = 8'h2;
                    16'h880B: data_out = 8'h3;
                    16'h880C: data_out = 8'h4;
                    16'h880D: data_out = 8'h5;
                    16'h880E: data_out = 8'h6;
                    16'h880F: data_out = 8'h7;
                    16'h8810: data_out = 8'h8;
                    16'h8811: data_out = 8'h9;
                    16'h8812: data_out = 8'hA;
                    16'h8813: data_out = 8'hB;
                    16'h8814: data_out = 8'hC;
                    16'h8815: data_out = 8'hD;
                    16'h8816: data_out = 8'hE;
                    16'h8817: data_out = 8'hF;
                    16'h8818: data_out = 8'h10;
                    16'h8819: data_out = 8'h11;
                    16'h881A: data_out = 8'h12;
                    16'h881B: data_out = 8'h13;
                    16'h881C: data_out = 8'h14;
                    16'h881D: data_out = 8'h15;
                    16'h881E: data_out = 8'h16;
                    16'h881F: data_out = 8'h17;
                    16'h8820: data_out = 8'h18;
                    16'h8821: data_out = 8'h19;
                    16'h8822: data_out = 8'h1A;
                    16'h8823: data_out = 8'h1B;
                    16'h8824: data_out = 8'h1C;
                    16'h8825: data_out = 8'h1D;
                    16'h8826: data_out = 8'h1E;
                    16'h8827: data_out = 8'h1F;
                    16'h8828: data_out = 8'h20;
                    16'h8829: data_out = 8'h21;
                    16'h882A: data_out = 8'h22;
                    16'h882B: data_out = 8'h23;
                    16'h882C: data_out = 8'h24;
                    16'h882D: data_out = 8'h25;
                    16'h882E: data_out = 8'h26;
                    16'h882F: data_out = 8'h27;
                    16'h8830: data_out = 8'h28;
                    16'h8831: data_out = 8'h29;
                    16'h8832: data_out = 8'h2A;
                    16'h8833: data_out = 8'h2B;
                    16'h8834: data_out = 8'h2C;
                    16'h8835: data_out = 8'h2D;
                    16'h8836: data_out = 8'h2E;
                    16'h8837: data_out = 8'h2F;
                    16'h8838: data_out = 8'h30;
                    16'h8839: data_out = 8'h31;
                    16'h883A: data_out = 8'h32;
                    16'h883B: data_out = 8'h33;
                    16'h883C: data_out = 8'h34;
                    16'h883D: data_out = 8'h35;
                    16'h883E: data_out = 8'h36;
                    16'h883F: data_out = 8'h37;
                    16'h8840: data_out = 8'h38;
                    16'h8841: data_out = 8'h39;
                    16'h8842: data_out = 8'h3A;
                    16'h8843: data_out = 8'h3B;
                    16'h8844: data_out = 8'h3C;
                    16'h8845: data_out = 8'h3D;
                    16'h8846: data_out = 8'h3E;
                    16'h8847: data_out = 8'h3F;
                    16'h8848: data_out = 8'h40;
                    16'h8849: data_out = 8'h41;
                    16'h884A: data_out = 8'h42;
                    16'h884B: data_out = 8'h43;
                    16'h884C: data_out = 8'h44;
                    16'h884D: data_out = 8'h45;
                    16'h884E: data_out = 8'h46;
                    16'h884F: data_out = 8'h47;
                    16'h8850: data_out = 8'h48;
                    16'h8851: data_out = 8'h49;
                    16'h8852: data_out = 8'h4A;
                    16'h8853: data_out = 8'h4B;
                    16'h8854: data_out = 8'h4C;
                    16'h8855: data_out = 8'h4D;
                    16'h8856: data_out = 8'h4E;
                    16'h8857: data_out = 8'h4F;
                    16'h8858: data_out = 8'h50;
                    16'h8859: data_out = 8'h51;
                    16'h885A: data_out = 8'h52;
                    16'h885B: data_out = 8'h53;
                    16'h885C: data_out = 8'h54;
                    16'h885D: data_out = 8'h55;
                    16'h885E: data_out = 8'h56;
                    16'h885F: data_out = 8'h57;
                    16'h8860: data_out = 8'h58;
                    16'h8861: data_out = 8'h59;
                    16'h8862: data_out = 8'h5A;
                    16'h8863: data_out = 8'h5B;
                    16'h8864: data_out = 8'h5C;
                    16'h8865: data_out = 8'h5D;
                    16'h8866: data_out = 8'h5E;
                    16'h8867: data_out = 8'h5F;
                    16'h8868: data_out = 8'h60;
                    16'h8869: data_out = 8'h61;
                    16'h886A: data_out = 8'h62;
                    16'h886B: data_out = 8'h63;
                    16'h886C: data_out = 8'h64;
                    16'h886D: data_out = 8'h65;
                    16'h886E: data_out = 8'h66;
                    16'h886F: data_out = 8'h67;
                    16'h8870: data_out = 8'h68;
                    16'h8871: data_out = 8'h69;
                    16'h8872: data_out = 8'h6A;
                    16'h8873: data_out = 8'h6B;
                    16'h8874: data_out = 8'h6C;
                    16'h8875: data_out = 8'h6D;
                    16'h8876: data_out = 8'h6E;
                    16'h8877: data_out = 8'h6F;
                    16'h8878: data_out = 8'h70;
                    16'h8879: data_out = 8'h71;
                    16'h887A: data_out = 8'h72;
                    16'h887B: data_out = 8'h73;
                    16'h887C: data_out = 8'h74;
                    16'h887D: data_out = 8'h75;
                    16'h887E: data_out = 8'h76;
                    16'h887F: data_out = 8'h77;
                    16'h8880: data_out = 8'h88;
                    16'h8881: data_out = 8'h89;
                    16'h8882: data_out = 8'h8A;
                    16'h8883: data_out = 8'h8B;
                    16'h8884: data_out = 8'h8C;
                    16'h8885: data_out = 8'h8D;
                    16'h8886: data_out = 8'h8E;
                    16'h8887: data_out = 8'h8F;
                    16'h8888: data_out = 8'h90;
                    16'h8889: data_out = 8'h91;
                    16'h888A: data_out = 8'h92;
                    16'h888B: data_out = 8'h93;
                    16'h888C: data_out = 8'h94;
                    16'h888D: data_out = 8'h95;
                    16'h888E: data_out = 8'h96;
                    16'h888F: data_out = 8'h97;
                    16'h8890: data_out = 8'h98;
                    16'h8891: data_out = 8'h99;
                    16'h8892: data_out = 8'h9A;
                    16'h8893: data_out = 8'h9B;
                    16'h8894: data_out = 8'h9C;
                    16'h8895: data_out = 8'h9D;
                    16'h8896: data_out = 8'h9E;
                    16'h8897: data_out = 8'h9F;
                    16'h8898: data_out = 8'hA0;
                    16'h8899: data_out = 8'hA1;
                    16'h889A: data_out = 8'hA2;
                    16'h889B: data_out = 8'hA3;
                    16'h889C: data_out = 8'hA4;
                    16'h889D: data_out = 8'hA5;
                    16'h889E: data_out = 8'hA6;
                    16'h889F: data_out = 8'hA7;
                    16'h88A0: data_out = 8'hA8;
                    16'h88A1: data_out = 8'hA9;
                    16'h88A2: data_out = 8'hAA;
                    16'h88A3: data_out = 8'hAB;
                    16'h88A4: data_out = 8'hAC;
                    16'h88A5: data_out = 8'hAD;
                    16'h88A6: data_out = 8'hAE;
                    16'h88A7: data_out = 8'hAF;
                    16'h88A8: data_out = 8'hB0;
                    16'h88A9: data_out = 8'hB1;
                    16'h88AA: data_out = 8'hB2;
                    16'h88AB: data_out = 8'hB3;
                    16'h88AC: data_out = 8'hB4;
                    16'h88AD: data_out = 8'hB5;
                    16'h88AE: data_out = 8'hB6;
                    16'h88AF: data_out = 8'hB7;
                    16'h88B0: data_out = 8'hB8;
                    16'h88B1: data_out = 8'hB9;
                    16'h88B2: data_out = 8'hBA;
                    16'h88B3: data_out = 8'hBB;
                    16'h88B4: data_out = 8'hBC;
                    16'h88B5: data_out = 8'hBD;
                    16'h88B6: data_out = 8'hBE;
                    16'h88B7: data_out = 8'hBF;
                    16'h88B8: data_out = 8'hC0;
                    16'h88B9: data_out = 8'hC1;
                    16'h88BA: data_out = 8'hC2;
                    16'h88BB: data_out = 8'hC3;
                    16'h88BC: data_out = 8'hC4;
                    16'h88BD: data_out = 8'hC5;
                    16'h88BE: data_out = 8'hC6;
                    16'h88BF: data_out = 8'hC7;
                    16'h88C0: data_out = 8'hC8;
                    16'h88C1: data_out = 8'hC9;
                    16'h88C2: data_out = 8'hCA;
                    16'h88C3: data_out = 8'hCB;
                    16'h88C4: data_out = 8'hCC;
                    16'h88C5: data_out = 8'hCD;
                    16'h88C6: data_out = 8'hCE;
                    16'h88C7: data_out = 8'hCF;
                    16'h88C8: data_out = 8'hD0;
                    16'h88C9: data_out = 8'hD1;
                    16'h88CA: data_out = 8'hD2;
                    16'h88CB: data_out = 8'hD3;
                    16'h88CC: data_out = 8'hD4;
                    16'h88CD: data_out = 8'hD5;
                    16'h88CE: data_out = 8'hD6;
                    16'h88CF: data_out = 8'hD7;
                    16'h88D0: data_out = 8'hD8;
                    16'h88D1: data_out = 8'hD9;
                    16'h88D2: data_out = 8'hDA;
                    16'h88D3: data_out = 8'hDB;
                    16'h88D4: data_out = 8'hDC;
                    16'h88D5: data_out = 8'hDD;
                    16'h88D6: data_out = 8'hDE;
                    16'h88D7: data_out = 8'hDF;
                    16'h88D8: data_out = 8'hE0;
                    16'h88D9: data_out = 8'hE1;
                    16'h88DA: data_out = 8'hE2;
                    16'h88DB: data_out = 8'hE3;
                    16'h88DC: data_out = 8'hE4;
                    16'h88DD: data_out = 8'hE5;
                    16'h88DE: data_out = 8'hE6;
                    16'h88DF: data_out = 8'hE7;
                    16'h88E0: data_out = 8'hE8;
                    16'h88E1: data_out = 8'hE9;
                    16'h88E2: data_out = 8'hEA;
                    16'h88E3: data_out = 8'hEB;
                    16'h88E4: data_out = 8'hEC;
                    16'h88E5: data_out = 8'hED;
                    16'h88E6: data_out = 8'hEE;
                    16'h88E7: data_out = 8'hEF;
                    16'h88E8: data_out = 8'hF0;
                    16'h88E9: data_out = 8'hF1;
                    16'h88EA: data_out = 8'hF2;
                    16'h88EB: data_out = 8'hF3;
                    16'h88EC: data_out = 8'hF4;
                    16'h88ED: data_out = 8'hF5;
                    16'h88EE: data_out = 8'hF6;
                    16'h88EF: data_out = 8'hF7;
                    16'h88F0: data_out = 8'hF8;
                    16'h88F1: data_out = 8'hF9;
                    16'h88F2: data_out = 8'hFA;
                    16'h88F3: data_out = 8'hFB;
                    16'h88F4: data_out = 8'hFC;
                    16'h88F5: data_out = 8'hFD;
                    16'h88F6: data_out = 8'hFE;
                    16'h88F7: data_out = 8'hFF;
                    16'h88F8: data_out = 8'h80;
                    16'h88F9: data_out = 8'h81;
                    16'h88FA: data_out = 8'h82;
                    16'h88FB: data_out = 8'h83;
                    16'h88FC: data_out = 8'h84;
                    16'h88FD: data_out = 8'h85;
                    16'h88FE: data_out = 8'h86;
                    16'h88FF: data_out = 8'h87;
                    16'h8900: data_out = 8'h89;
                    16'h8901: data_out = 8'h88;
                    16'h8902: data_out = 8'h87;
                    16'h8903: data_out = 8'h86;
                    16'h8904: data_out = 8'h85;
                    16'h8905: data_out = 8'h84;
                    16'h8906: data_out = 8'h83;
                    16'h8907: data_out = 8'h82;
                    16'h8908: data_out = 8'h81;
                    16'h8909: data_out = 8'h0;
                    16'h890A: data_out = 8'h1;
                    16'h890B: data_out = 8'h2;
                    16'h890C: data_out = 8'h3;
                    16'h890D: data_out = 8'h4;
                    16'h890E: data_out = 8'h5;
                    16'h890F: data_out = 8'h6;
                    16'h8910: data_out = 8'h7;
                    16'h8911: data_out = 8'h8;
                    16'h8912: data_out = 8'h9;
                    16'h8913: data_out = 8'hA;
                    16'h8914: data_out = 8'hB;
                    16'h8915: data_out = 8'hC;
                    16'h8916: data_out = 8'hD;
                    16'h8917: data_out = 8'hE;
                    16'h8918: data_out = 8'hF;
                    16'h8919: data_out = 8'h10;
                    16'h891A: data_out = 8'h11;
                    16'h891B: data_out = 8'h12;
                    16'h891C: data_out = 8'h13;
                    16'h891D: data_out = 8'h14;
                    16'h891E: data_out = 8'h15;
                    16'h891F: data_out = 8'h16;
                    16'h8920: data_out = 8'h17;
                    16'h8921: data_out = 8'h18;
                    16'h8922: data_out = 8'h19;
                    16'h8923: data_out = 8'h1A;
                    16'h8924: data_out = 8'h1B;
                    16'h8925: data_out = 8'h1C;
                    16'h8926: data_out = 8'h1D;
                    16'h8927: data_out = 8'h1E;
                    16'h8928: data_out = 8'h1F;
                    16'h8929: data_out = 8'h20;
                    16'h892A: data_out = 8'h21;
                    16'h892B: data_out = 8'h22;
                    16'h892C: data_out = 8'h23;
                    16'h892D: data_out = 8'h24;
                    16'h892E: data_out = 8'h25;
                    16'h892F: data_out = 8'h26;
                    16'h8930: data_out = 8'h27;
                    16'h8931: data_out = 8'h28;
                    16'h8932: data_out = 8'h29;
                    16'h8933: data_out = 8'h2A;
                    16'h8934: data_out = 8'h2B;
                    16'h8935: data_out = 8'h2C;
                    16'h8936: data_out = 8'h2D;
                    16'h8937: data_out = 8'h2E;
                    16'h8938: data_out = 8'h2F;
                    16'h8939: data_out = 8'h30;
                    16'h893A: data_out = 8'h31;
                    16'h893B: data_out = 8'h32;
                    16'h893C: data_out = 8'h33;
                    16'h893D: data_out = 8'h34;
                    16'h893E: data_out = 8'h35;
                    16'h893F: data_out = 8'h36;
                    16'h8940: data_out = 8'h37;
                    16'h8941: data_out = 8'h38;
                    16'h8942: data_out = 8'h39;
                    16'h8943: data_out = 8'h3A;
                    16'h8944: data_out = 8'h3B;
                    16'h8945: data_out = 8'h3C;
                    16'h8946: data_out = 8'h3D;
                    16'h8947: data_out = 8'h3E;
                    16'h8948: data_out = 8'h3F;
                    16'h8949: data_out = 8'h40;
                    16'h894A: data_out = 8'h41;
                    16'h894B: data_out = 8'h42;
                    16'h894C: data_out = 8'h43;
                    16'h894D: data_out = 8'h44;
                    16'h894E: data_out = 8'h45;
                    16'h894F: data_out = 8'h46;
                    16'h8950: data_out = 8'h47;
                    16'h8951: data_out = 8'h48;
                    16'h8952: data_out = 8'h49;
                    16'h8953: data_out = 8'h4A;
                    16'h8954: data_out = 8'h4B;
                    16'h8955: data_out = 8'h4C;
                    16'h8956: data_out = 8'h4D;
                    16'h8957: data_out = 8'h4E;
                    16'h8958: data_out = 8'h4F;
                    16'h8959: data_out = 8'h50;
                    16'h895A: data_out = 8'h51;
                    16'h895B: data_out = 8'h52;
                    16'h895C: data_out = 8'h53;
                    16'h895D: data_out = 8'h54;
                    16'h895E: data_out = 8'h55;
                    16'h895F: data_out = 8'h56;
                    16'h8960: data_out = 8'h57;
                    16'h8961: data_out = 8'h58;
                    16'h8962: data_out = 8'h59;
                    16'h8963: data_out = 8'h5A;
                    16'h8964: data_out = 8'h5B;
                    16'h8965: data_out = 8'h5C;
                    16'h8966: data_out = 8'h5D;
                    16'h8967: data_out = 8'h5E;
                    16'h8968: data_out = 8'h5F;
                    16'h8969: data_out = 8'h60;
                    16'h896A: data_out = 8'h61;
                    16'h896B: data_out = 8'h62;
                    16'h896C: data_out = 8'h63;
                    16'h896D: data_out = 8'h64;
                    16'h896E: data_out = 8'h65;
                    16'h896F: data_out = 8'h66;
                    16'h8970: data_out = 8'h67;
                    16'h8971: data_out = 8'h68;
                    16'h8972: data_out = 8'h69;
                    16'h8973: data_out = 8'h6A;
                    16'h8974: data_out = 8'h6B;
                    16'h8975: data_out = 8'h6C;
                    16'h8976: data_out = 8'h6D;
                    16'h8977: data_out = 8'h6E;
                    16'h8978: data_out = 8'h6F;
                    16'h8979: data_out = 8'h70;
                    16'h897A: data_out = 8'h71;
                    16'h897B: data_out = 8'h72;
                    16'h897C: data_out = 8'h73;
                    16'h897D: data_out = 8'h74;
                    16'h897E: data_out = 8'h75;
                    16'h897F: data_out = 8'h76;
                    16'h8980: data_out = 8'h89;
                    16'h8981: data_out = 8'h8A;
                    16'h8982: data_out = 8'h8B;
                    16'h8983: data_out = 8'h8C;
                    16'h8984: data_out = 8'h8D;
                    16'h8985: data_out = 8'h8E;
                    16'h8986: data_out = 8'h8F;
                    16'h8987: data_out = 8'h90;
                    16'h8988: data_out = 8'h91;
                    16'h8989: data_out = 8'h92;
                    16'h898A: data_out = 8'h93;
                    16'h898B: data_out = 8'h94;
                    16'h898C: data_out = 8'h95;
                    16'h898D: data_out = 8'h96;
                    16'h898E: data_out = 8'h97;
                    16'h898F: data_out = 8'h98;
                    16'h8990: data_out = 8'h99;
                    16'h8991: data_out = 8'h9A;
                    16'h8992: data_out = 8'h9B;
                    16'h8993: data_out = 8'h9C;
                    16'h8994: data_out = 8'h9D;
                    16'h8995: data_out = 8'h9E;
                    16'h8996: data_out = 8'h9F;
                    16'h8997: data_out = 8'hA0;
                    16'h8998: data_out = 8'hA1;
                    16'h8999: data_out = 8'hA2;
                    16'h899A: data_out = 8'hA3;
                    16'h899B: data_out = 8'hA4;
                    16'h899C: data_out = 8'hA5;
                    16'h899D: data_out = 8'hA6;
                    16'h899E: data_out = 8'hA7;
                    16'h899F: data_out = 8'hA8;
                    16'h89A0: data_out = 8'hA9;
                    16'h89A1: data_out = 8'hAA;
                    16'h89A2: data_out = 8'hAB;
                    16'h89A3: data_out = 8'hAC;
                    16'h89A4: data_out = 8'hAD;
                    16'h89A5: data_out = 8'hAE;
                    16'h89A6: data_out = 8'hAF;
                    16'h89A7: data_out = 8'hB0;
                    16'h89A8: data_out = 8'hB1;
                    16'h89A9: data_out = 8'hB2;
                    16'h89AA: data_out = 8'hB3;
                    16'h89AB: data_out = 8'hB4;
                    16'h89AC: data_out = 8'hB5;
                    16'h89AD: data_out = 8'hB6;
                    16'h89AE: data_out = 8'hB7;
                    16'h89AF: data_out = 8'hB8;
                    16'h89B0: data_out = 8'hB9;
                    16'h89B1: data_out = 8'hBA;
                    16'h89B2: data_out = 8'hBB;
                    16'h89B3: data_out = 8'hBC;
                    16'h89B4: data_out = 8'hBD;
                    16'h89B5: data_out = 8'hBE;
                    16'h89B6: data_out = 8'hBF;
                    16'h89B7: data_out = 8'hC0;
                    16'h89B8: data_out = 8'hC1;
                    16'h89B9: data_out = 8'hC2;
                    16'h89BA: data_out = 8'hC3;
                    16'h89BB: data_out = 8'hC4;
                    16'h89BC: data_out = 8'hC5;
                    16'h89BD: data_out = 8'hC6;
                    16'h89BE: data_out = 8'hC7;
                    16'h89BF: data_out = 8'hC8;
                    16'h89C0: data_out = 8'hC9;
                    16'h89C1: data_out = 8'hCA;
                    16'h89C2: data_out = 8'hCB;
                    16'h89C3: data_out = 8'hCC;
                    16'h89C4: data_out = 8'hCD;
                    16'h89C5: data_out = 8'hCE;
                    16'h89C6: data_out = 8'hCF;
                    16'h89C7: data_out = 8'hD0;
                    16'h89C8: data_out = 8'hD1;
                    16'h89C9: data_out = 8'hD2;
                    16'h89CA: data_out = 8'hD3;
                    16'h89CB: data_out = 8'hD4;
                    16'h89CC: data_out = 8'hD5;
                    16'h89CD: data_out = 8'hD6;
                    16'h89CE: data_out = 8'hD7;
                    16'h89CF: data_out = 8'hD8;
                    16'h89D0: data_out = 8'hD9;
                    16'h89D1: data_out = 8'hDA;
                    16'h89D2: data_out = 8'hDB;
                    16'h89D3: data_out = 8'hDC;
                    16'h89D4: data_out = 8'hDD;
                    16'h89D5: data_out = 8'hDE;
                    16'h89D6: data_out = 8'hDF;
                    16'h89D7: data_out = 8'hE0;
                    16'h89D8: data_out = 8'hE1;
                    16'h89D9: data_out = 8'hE2;
                    16'h89DA: data_out = 8'hE3;
                    16'h89DB: data_out = 8'hE4;
                    16'h89DC: data_out = 8'hE5;
                    16'h89DD: data_out = 8'hE6;
                    16'h89DE: data_out = 8'hE7;
                    16'h89DF: data_out = 8'hE8;
                    16'h89E0: data_out = 8'hE9;
                    16'h89E1: data_out = 8'hEA;
                    16'h89E2: data_out = 8'hEB;
                    16'h89E3: data_out = 8'hEC;
                    16'h89E4: data_out = 8'hED;
                    16'h89E5: data_out = 8'hEE;
                    16'h89E6: data_out = 8'hEF;
                    16'h89E7: data_out = 8'hF0;
                    16'h89E8: data_out = 8'hF1;
                    16'h89E9: data_out = 8'hF2;
                    16'h89EA: data_out = 8'hF3;
                    16'h89EB: data_out = 8'hF4;
                    16'h89EC: data_out = 8'hF5;
                    16'h89ED: data_out = 8'hF6;
                    16'h89EE: data_out = 8'hF7;
                    16'h89EF: data_out = 8'hF8;
                    16'h89F0: data_out = 8'hF9;
                    16'h89F1: data_out = 8'hFA;
                    16'h89F2: data_out = 8'hFB;
                    16'h89F3: data_out = 8'hFC;
                    16'h89F4: data_out = 8'hFD;
                    16'h89F5: data_out = 8'hFE;
                    16'h89F6: data_out = 8'hFF;
                    16'h89F7: data_out = 8'h80;
                    16'h89F8: data_out = 8'h81;
                    16'h89F9: data_out = 8'h82;
                    16'h89FA: data_out = 8'h83;
                    16'h89FB: data_out = 8'h84;
                    16'h89FC: data_out = 8'h85;
                    16'h89FD: data_out = 8'h86;
                    16'h89FE: data_out = 8'h87;
                    16'h89FF: data_out = 8'h88;
                    16'h8A00: data_out = 8'h8A;
                    16'h8A01: data_out = 8'h89;
                    16'h8A02: data_out = 8'h88;
                    16'h8A03: data_out = 8'h87;
                    16'h8A04: data_out = 8'h86;
                    16'h8A05: data_out = 8'h85;
                    16'h8A06: data_out = 8'h84;
                    16'h8A07: data_out = 8'h83;
                    16'h8A08: data_out = 8'h82;
                    16'h8A09: data_out = 8'h81;
                    16'h8A0A: data_out = 8'h0;
                    16'h8A0B: data_out = 8'h1;
                    16'h8A0C: data_out = 8'h2;
                    16'h8A0D: data_out = 8'h3;
                    16'h8A0E: data_out = 8'h4;
                    16'h8A0F: data_out = 8'h5;
                    16'h8A10: data_out = 8'h6;
                    16'h8A11: data_out = 8'h7;
                    16'h8A12: data_out = 8'h8;
                    16'h8A13: data_out = 8'h9;
                    16'h8A14: data_out = 8'hA;
                    16'h8A15: data_out = 8'hB;
                    16'h8A16: data_out = 8'hC;
                    16'h8A17: data_out = 8'hD;
                    16'h8A18: data_out = 8'hE;
                    16'h8A19: data_out = 8'hF;
                    16'h8A1A: data_out = 8'h10;
                    16'h8A1B: data_out = 8'h11;
                    16'h8A1C: data_out = 8'h12;
                    16'h8A1D: data_out = 8'h13;
                    16'h8A1E: data_out = 8'h14;
                    16'h8A1F: data_out = 8'h15;
                    16'h8A20: data_out = 8'h16;
                    16'h8A21: data_out = 8'h17;
                    16'h8A22: data_out = 8'h18;
                    16'h8A23: data_out = 8'h19;
                    16'h8A24: data_out = 8'h1A;
                    16'h8A25: data_out = 8'h1B;
                    16'h8A26: data_out = 8'h1C;
                    16'h8A27: data_out = 8'h1D;
                    16'h8A28: data_out = 8'h1E;
                    16'h8A29: data_out = 8'h1F;
                    16'h8A2A: data_out = 8'h20;
                    16'h8A2B: data_out = 8'h21;
                    16'h8A2C: data_out = 8'h22;
                    16'h8A2D: data_out = 8'h23;
                    16'h8A2E: data_out = 8'h24;
                    16'h8A2F: data_out = 8'h25;
                    16'h8A30: data_out = 8'h26;
                    16'h8A31: data_out = 8'h27;
                    16'h8A32: data_out = 8'h28;
                    16'h8A33: data_out = 8'h29;
                    16'h8A34: data_out = 8'h2A;
                    16'h8A35: data_out = 8'h2B;
                    16'h8A36: data_out = 8'h2C;
                    16'h8A37: data_out = 8'h2D;
                    16'h8A38: data_out = 8'h2E;
                    16'h8A39: data_out = 8'h2F;
                    16'h8A3A: data_out = 8'h30;
                    16'h8A3B: data_out = 8'h31;
                    16'h8A3C: data_out = 8'h32;
                    16'h8A3D: data_out = 8'h33;
                    16'h8A3E: data_out = 8'h34;
                    16'h8A3F: data_out = 8'h35;
                    16'h8A40: data_out = 8'h36;
                    16'h8A41: data_out = 8'h37;
                    16'h8A42: data_out = 8'h38;
                    16'h8A43: data_out = 8'h39;
                    16'h8A44: data_out = 8'h3A;
                    16'h8A45: data_out = 8'h3B;
                    16'h8A46: data_out = 8'h3C;
                    16'h8A47: data_out = 8'h3D;
                    16'h8A48: data_out = 8'h3E;
                    16'h8A49: data_out = 8'h3F;
                    16'h8A4A: data_out = 8'h40;
                    16'h8A4B: data_out = 8'h41;
                    16'h8A4C: data_out = 8'h42;
                    16'h8A4D: data_out = 8'h43;
                    16'h8A4E: data_out = 8'h44;
                    16'h8A4F: data_out = 8'h45;
                    16'h8A50: data_out = 8'h46;
                    16'h8A51: data_out = 8'h47;
                    16'h8A52: data_out = 8'h48;
                    16'h8A53: data_out = 8'h49;
                    16'h8A54: data_out = 8'h4A;
                    16'h8A55: data_out = 8'h4B;
                    16'h8A56: data_out = 8'h4C;
                    16'h8A57: data_out = 8'h4D;
                    16'h8A58: data_out = 8'h4E;
                    16'h8A59: data_out = 8'h4F;
                    16'h8A5A: data_out = 8'h50;
                    16'h8A5B: data_out = 8'h51;
                    16'h8A5C: data_out = 8'h52;
                    16'h8A5D: data_out = 8'h53;
                    16'h8A5E: data_out = 8'h54;
                    16'h8A5F: data_out = 8'h55;
                    16'h8A60: data_out = 8'h56;
                    16'h8A61: data_out = 8'h57;
                    16'h8A62: data_out = 8'h58;
                    16'h8A63: data_out = 8'h59;
                    16'h8A64: data_out = 8'h5A;
                    16'h8A65: data_out = 8'h5B;
                    16'h8A66: data_out = 8'h5C;
                    16'h8A67: data_out = 8'h5D;
                    16'h8A68: data_out = 8'h5E;
                    16'h8A69: data_out = 8'h5F;
                    16'h8A6A: data_out = 8'h60;
                    16'h8A6B: data_out = 8'h61;
                    16'h8A6C: data_out = 8'h62;
                    16'h8A6D: data_out = 8'h63;
                    16'h8A6E: data_out = 8'h64;
                    16'h8A6F: data_out = 8'h65;
                    16'h8A70: data_out = 8'h66;
                    16'h8A71: data_out = 8'h67;
                    16'h8A72: data_out = 8'h68;
                    16'h8A73: data_out = 8'h69;
                    16'h8A74: data_out = 8'h6A;
                    16'h8A75: data_out = 8'h6B;
                    16'h8A76: data_out = 8'h6C;
                    16'h8A77: data_out = 8'h6D;
                    16'h8A78: data_out = 8'h6E;
                    16'h8A79: data_out = 8'h6F;
                    16'h8A7A: data_out = 8'h70;
                    16'h8A7B: data_out = 8'h71;
                    16'h8A7C: data_out = 8'h72;
                    16'h8A7D: data_out = 8'h73;
                    16'h8A7E: data_out = 8'h74;
                    16'h8A7F: data_out = 8'h75;
                    16'h8A80: data_out = 8'h8A;
                    16'h8A81: data_out = 8'h8B;
                    16'h8A82: data_out = 8'h8C;
                    16'h8A83: data_out = 8'h8D;
                    16'h8A84: data_out = 8'h8E;
                    16'h8A85: data_out = 8'h8F;
                    16'h8A86: data_out = 8'h90;
                    16'h8A87: data_out = 8'h91;
                    16'h8A88: data_out = 8'h92;
                    16'h8A89: data_out = 8'h93;
                    16'h8A8A: data_out = 8'h94;
                    16'h8A8B: data_out = 8'h95;
                    16'h8A8C: data_out = 8'h96;
                    16'h8A8D: data_out = 8'h97;
                    16'h8A8E: data_out = 8'h98;
                    16'h8A8F: data_out = 8'h99;
                    16'h8A90: data_out = 8'h9A;
                    16'h8A91: data_out = 8'h9B;
                    16'h8A92: data_out = 8'h9C;
                    16'h8A93: data_out = 8'h9D;
                    16'h8A94: data_out = 8'h9E;
                    16'h8A95: data_out = 8'h9F;
                    16'h8A96: data_out = 8'hA0;
                    16'h8A97: data_out = 8'hA1;
                    16'h8A98: data_out = 8'hA2;
                    16'h8A99: data_out = 8'hA3;
                    16'h8A9A: data_out = 8'hA4;
                    16'h8A9B: data_out = 8'hA5;
                    16'h8A9C: data_out = 8'hA6;
                    16'h8A9D: data_out = 8'hA7;
                    16'h8A9E: data_out = 8'hA8;
                    16'h8A9F: data_out = 8'hA9;
                    16'h8AA0: data_out = 8'hAA;
                    16'h8AA1: data_out = 8'hAB;
                    16'h8AA2: data_out = 8'hAC;
                    16'h8AA3: data_out = 8'hAD;
                    16'h8AA4: data_out = 8'hAE;
                    16'h8AA5: data_out = 8'hAF;
                    16'h8AA6: data_out = 8'hB0;
                    16'h8AA7: data_out = 8'hB1;
                    16'h8AA8: data_out = 8'hB2;
                    16'h8AA9: data_out = 8'hB3;
                    16'h8AAA: data_out = 8'hB4;
                    16'h8AAB: data_out = 8'hB5;
                    16'h8AAC: data_out = 8'hB6;
                    16'h8AAD: data_out = 8'hB7;
                    16'h8AAE: data_out = 8'hB8;
                    16'h8AAF: data_out = 8'hB9;
                    16'h8AB0: data_out = 8'hBA;
                    16'h8AB1: data_out = 8'hBB;
                    16'h8AB2: data_out = 8'hBC;
                    16'h8AB3: data_out = 8'hBD;
                    16'h8AB4: data_out = 8'hBE;
                    16'h8AB5: data_out = 8'hBF;
                    16'h8AB6: data_out = 8'hC0;
                    16'h8AB7: data_out = 8'hC1;
                    16'h8AB8: data_out = 8'hC2;
                    16'h8AB9: data_out = 8'hC3;
                    16'h8ABA: data_out = 8'hC4;
                    16'h8ABB: data_out = 8'hC5;
                    16'h8ABC: data_out = 8'hC6;
                    16'h8ABD: data_out = 8'hC7;
                    16'h8ABE: data_out = 8'hC8;
                    16'h8ABF: data_out = 8'hC9;
                    16'h8AC0: data_out = 8'hCA;
                    16'h8AC1: data_out = 8'hCB;
                    16'h8AC2: data_out = 8'hCC;
                    16'h8AC3: data_out = 8'hCD;
                    16'h8AC4: data_out = 8'hCE;
                    16'h8AC5: data_out = 8'hCF;
                    16'h8AC6: data_out = 8'hD0;
                    16'h8AC7: data_out = 8'hD1;
                    16'h8AC8: data_out = 8'hD2;
                    16'h8AC9: data_out = 8'hD3;
                    16'h8ACA: data_out = 8'hD4;
                    16'h8ACB: data_out = 8'hD5;
                    16'h8ACC: data_out = 8'hD6;
                    16'h8ACD: data_out = 8'hD7;
                    16'h8ACE: data_out = 8'hD8;
                    16'h8ACF: data_out = 8'hD9;
                    16'h8AD0: data_out = 8'hDA;
                    16'h8AD1: data_out = 8'hDB;
                    16'h8AD2: data_out = 8'hDC;
                    16'h8AD3: data_out = 8'hDD;
                    16'h8AD4: data_out = 8'hDE;
                    16'h8AD5: data_out = 8'hDF;
                    16'h8AD6: data_out = 8'hE0;
                    16'h8AD7: data_out = 8'hE1;
                    16'h8AD8: data_out = 8'hE2;
                    16'h8AD9: data_out = 8'hE3;
                    16'h8ADA: data_out = 8'hE4;
                    16'h8ADB: data_out = 8'hE5;
                    16'h8ADC: data_out = 8'hE6;
                    16'h8ADD: data_out = 8'hE7;
                    16'h8ADE: data_out = 8'hE8;
                    16'h8ADF: data_out = 8'hE9;
                    16'h8AE0: data_out = 8'hEA;
                    16'h8AE1: data_out = 8'hEB;
                    16'h8AE2: data_out = 8'hEC;
                    16'h8AE3: data_out = 8'hED;
                    16'h8AE4: data_out = 8'hEE;
                    16'h8AE5: data_out = 8'hEF;
                    16'h8AE6: data_out = 8'hF0;
                    16'h8AE7: data_out = 8'hF1;
                    16'h8AE8: data_out = 8'hF2;
                    16'h8AE9: data_out = 8'hF3;
                    16'h8AEA: data_out = 8'hF4;
                    16'h8AEB: data_out = 8'hF5;
                    16'h8AEC: data_out = 8'hF6;
                    16'h8AED: data_out = 8'hF7;
                    16'h8AEE: data_out = 8'hF8;
                    16'h8AEF: data_out = 8'hF9;
                    16'h8AF0: data_out = 8'hFA;
                    16'h8AF1: data_out = 8'hFB;
                    16'h8AF2: data_out = 8'hFC;
                    16'h8AF3: data_out = 8'hFD;
                    16'h8AF4: data_out = 8'hFE;
                    16'h8AF5: data_out = 8'hFF;
                    16'h8AF6: data_out = 8'h80;
                    16'h8AF7: data_out = 8'h81;
                    16'h8AF8: data_out = 8'h82;
                    16'h8AF9: data_out = 8'h83;
                    16'h8AFA: data_out = 8'h84;
                    16'h8AFB: data_out = 8'h85;
                    16'h8AFC: data_out = 8'h86;
                    16'h8AFD: data_out = 8'h87;
                    16'h8AFE: data_out = 8'h88;
                    16'h8AFF: data_out = 8'h89;
                    16'h8B00: data_out = 8'h8B;
                    16'h8B01: data_out = 8'h8A;
                    16'h8B02: data_out = 8'h89;
                    16'h8B03: data_out = 8'h88;
                    16'h8B04: data_out = 8'h87;
                    16'h8B05: data_out = 8'h86;
                    16'h8B06: data_out = 8'h85;
                    16'h8B07: data_out = 8'h84;
                    16'h8B08: data_out = 8'h83;
                    16'h8B09: data_out = 8'h82;
                    16'h8B0A: data_out = 8'h81;
                    16'h8B0B: data_out = 8'h0;
                    16'h8B0C: data_out = 8'h1;
                    16'h8B0D: data_out = 8'h2;
                    16'h8B0E: data_out = 8'h3;
                    16'h8B0F: data_out = 8'h4;
                    16'h8B10: data_out = 8'h5;
                    16'h8B11: data_out = 8'h6;
                    16'h8B12: data_out = 8'h7;
                    16'h8B13: data_out = 8'h8;
                    16'h8B14: data_out = 8'h9;
                    16'h8B15: data_out = 8'hA;
                    16'h8B16: data_out = 8'hB;
                    16'h8B17: data_out = 8'hC;
                    16'h8B18: data_out = 8'hD;
                    16'h8B19: data_out = 8'hE;
                    16'h8B1A: data_out = 8'hF;
                    16'h8B1B: data_out = 8'h10;
                    16'h8B1C: data_out = 8'h11;
                    16'h8B1D: data_out = 8'h12;
                    16'h8B1E: data_out = 8'h13;
                    16'h8B1F: data_out = 8'h14;
                    16'h8B20: data_out = 8'h15;
                    16'h8B21: data_out = 8'h16;
                    16'h8B22: data_out = 8'h17;
                    16'h8B23: data_out = 8'h18;
                    16'h8B24: data_out = 8'h19;
                    16'h8B25: data_out = 8'h1A;
                    16'h8B26: data_out = 8'h1B;
                    16'h8B27: data_out = 8'h1C;
                    16'h8B28: data_out = 8'h1D;
                    16'h8B29: data_out = 8'h1E;
                    16'h8B2A: data_out = 8'h1F;
                    16'h8B2B: data_out = 8'h20;
                    16'h8B2C: data_out = 8'h21;
                    16'h8B2D: data_out = 8'h22;
                    16'h8B2E: data_out = 8'h23;
                    16'h8B2F: data_out = 8'h24;
                    16'h8B30: data_out = 8'h25;
                    16'h8B31: data_out = 8'h26;
                    16'h8B32: data_out = 8'h27;
                    16'h8B33: data_out = 8'h28;
                    16'h8B34: data_out = 8'h29;
                    16'h8B35: data_out = 8'h2A;
                    16'h8B36: data_out = 8'h2B;
                    16'h8B37: data_out = 8'h2C;
                    16'h8B38: data_out = 8'h2D;
                    16'h8B39: data_out = 8'h2E;
                    16'h8B3A: data_out = 8'h2F;
                    16'h8B3B: data_out = 8'h30;
                    16'h8B3C: data_out = 8'h31;
                    16'h8B3D: data_out = 8'h32;
                    16'h8B3E: data_out = 8'h33;
                    16'h8B3F: data_out = 8'h34;
                    16'h8B40: data_out = 8'h35;
                    16'h8B41: data_out = 8'h36;
                    16'h8B42: data_out = 8'h37;
                    16'h8B43: data_out = 8'h38;
                    16'h8B44: data_out = 8'h39;
                    16'h8B45: data_out = 8'h3A;
                    16'h8B46: data_out = 8'h3B;
                    16'h8B47: data_out = 8'h3C;
                    16'h8B48: data_out = 8'h3D;
                    16'h8B49: data_out = 8'h3E;
                    16'h8B4A: data_out = 8'h3F;
                    16'h8B4B: data_out = 8'h40;
                    16'h8B4C: data_out = 8'h41;
                    16'h8B4D: data_out = 8'h42;
                    16'h8B4E: data_out = 8'h43;
                    16'h8B4F: data_out = 8'h44;
                    16'h8B50: data_out = 8'h45;
                    16'h8B51: data_out = 8'h46;
                    16'h8B52: data_out = 8'h47;
                    16'h8B53: data_out = 8'h48;
                    16'h8B54: data_out = 8'h49;
                    16'h8B55: data_out = 8'h4A;
                    16'h8B56: data_out = 8'h4B;
                    16'h8B57: data_out = 8'h4C;
                    16'h8B58: data_out = 8'h4D;
                    16'h8B59: data_out = 8'h4E;
                    16'h8B5A: data_out = 8'h4F;
                    16'h8B5B: data_out = 8'h50;
                    16'h8B5C: data_out = 8'h51;
                    16'h8B5D: data_out = 8'h52;
                    16'h8B5E: data_out = 8'h53;
                    16'h8B5F: data_out = 8'h54;
                    16'h8B60: data_out = 8'h55;
                    16'h8B61: data_out = 8'h56;
                    16'h8B62: data_out = 8'h57;
                    16'h8B63: data_out = 8'h58;
                    16'h8B64: data_out = 8'h59;
                    16'h8B65: data_out = 8'h5A;
                    16'h8B66: data_out = 8'h5B;
                    16'h8B67: data_out = 8'h5C;
                    16'h8B68: data_out = 8'h5D;
                    16'h8B69: data_out = 8'h5E;
                    16'h8B6A: data_out = 8'h5F;
                    16'h8B6B: data_out = 8'h60;
                    16'h8B6C: data_out = 8'h61;
                    16'h8B6D: data_out = 8'h62;
                    16'h8B6E: data_out = 8'h63;
                    16'h8B6F: data_out = 8'h64;
                    16'h8B70: data_out = 8'h65;
                    16'h8B71: data_out = 8'h66;
                    16'h8B72: data_out = 8'h67;
                    16'h8B73: data_out = 8'h68;
                    16'h8B74: data_out = 8'h69;
                    16'h8B75: data_out = 8'h6A;
                    16'h8B76: data_out = 8'h6B;
                    16'h8B77: data_out = 8'h6C;
                    16'h8B78: data_out = 8'h6D;
                    16'h8B79: data_out = 8'h6E;
                    16'h8B7A: data_out = 8'h6F;
                    16'h8B7B: data_out = 8'h70;
                    16'h8B7C: data_out = 8'h71;
                    16'h8B7D: data_out = 8'h72;
                    16'h8B7E: data_out = 8'h73;
                    16'h8B7F: data_out = 8'h74;
                    16'h8B80: data_out = 8'h8B;
                    16'h8B81: data_out = 8'h8C;
                    16'h8B82: data_out = 8'h8D;
                    16'h8B83: data_out = 8'h8E;
                    16'h8B84: data_out = 8'h8F;
                    16'h8B85: data_out = 8'h90;
                    16'h8B86: data_out = 8'h91;
                    16'h8B87: data_out = 8'h92;
                    16'h8B88: data_out = 8'h93;
                    16'h8B89: data_out = 8'h94;
                    16'h8B8A: data_out = 8'h95;
                    16'h8B8B: data_out = 8'h96;
                    16'h8B8C: data_out = 8'h97;
                    16'h8B8D: data_out = 8'h98;
                    16'h8B8E: data_out = 8'h99;
                    16'h8B8F: data_out = 8'h9A;
                    16'h8B90: data_out = 8'h9B;
                    16'h8B91: data_out = 8'h9C;
                    16'h8B92: data_out = 8'h9D;
                    16'h8B93: data_out = 8'h9E;
                    16'h8B94: data_out = 8'h9F;
                    16'h8B95: data_out = 8'hA0;
                    16'h8B96: data_out = 8'hA1;
                    16'h8B97: data_out = 8'hA2;
                    16'h8B98: data_out = 8'hA3;
                    16'h8B99: data_out = 8'hA4;
                    16'h8B9A: data_out = 8'hA5;
                    16'h8B9B: data_out = 8'hA6;
                    16'h8B9C: data_out = 8'hA7;
                    16'h8B9D: data_out = 8'hA8;
                    16'h8B9E: data_out = 8'hA9;
                    16'h8B9F: data_out = 8'hAA;
                    16'h8BA0: data_out = 8'hAB;
                    16'h8BA1: data_out = 8'hAC;
                    16'h8BA2: data_out = 8'hAD;
                    16'h8BA3: data_out = 8'hAE;
                    16'h8BA4: data_out = 8'hAF;
                    16'h8BA5: data_out = 8'hB0;
                    16'h8BA6: data_out = 8'hB1;
                    16'h8BA7: data_out = 8'hB2;
                    16'h8BA8: data_out = 8'hB3;
                    16'h8BA9: data_out = 8'hB4;
                    16'h8BAA: data_out = 8'hB5;
                    16'h8BAB: data_out = 8'hB6;
                    16'h8BAC: data_out = 8'hB7;
                    16'h8BAD: data_out = 8'hB8;
                    16'h8BAE: data_out = 8'hB9;
                    16'h8BAF: data_out = 8'hBA;
                    16'h8BB0: data_out = 8'hBB;
                    16'h8BB1: data_out = 8'hBC;
                    16'h8BB2: data_out = 8'hBD;
                    16'h8BB3: data_out = 8'hBE;
                    16'h8BB4: data_out = 8'hBF;
                    16'h8BB5: data_out = 8'hC0;
                    16'h8BB6: data_out = 8'hC1;
                    16'h8BB7: data_out = 8'hC2;
                    16'h8BB8: data_out = 8'hC3;
                    16'h8BB9: data_out = 8'hC4;
                    16'h8BBA: data_out = 8'hC5;
                    16'h8BBB: data_out = 8'hC6;
                    16'h8BBC: data_out = 8'hC7;
                    16'h8BBD: data_out = 8'hC8;
                    16'h8BBE: data_out = 8'hC9;
                    16'h8BBF: data_out = 8'hCA;
                    16'h8BC0: data_out = 8'hCB;
                    16'h8BC1: data_out = 8'hCC;
                    16'h8BC2: data_out = 8'hCD;
                    16'h8BC3: data_out = 8'hCE;
                    16'h8BC4: data_out = 8'hCF;
                    16'h8BC5: data_out = 8'hD0;
                    16'h8BC6: data_out = 8'hD1;
                    16'h8BC7: data_out = 8'hD2;
                    16'h8BC8: data_out = 8'hD3;
                    16'h8BC9: data_out = 8'hD4;
                    16'h8BCA: data_out = 8'hD5;
                    16'h8BCB: data_out = 8'hD6;
                    16'h8BCC: data_out = 8'hD7;
                    16'h8BCD: data_out = 8'hD8;
                    16'h8BCE: data_out = 8'hD9;
                    16'h8BCF: data_out = 8'hDA;
                    16'h8BD0: data_out = 8'hDB;
                    16'h8BD1: data_out = 8'hDC;
                    16'h8BD2: data_out = 8'hDD;
                    16'h8BD3: data_out = 8'hDE;
                    16'h8BD4: data_out = 8'hDF;
                    16'h8BD5: data_out = 8'hE0;
                    16'h8BD6: data_out = 8'hE1;
                    16'h8BD7: data_out = 8'hE2;
                    16'h8BD8: data_out = 8'hE3;
                    16'h8BD9: data_out = 8'hE4;
                    16'h8BDA: data_out = 8'hE5;
                    16'h8BDB: data_out = 8'hE6;
                    16'h8BDC: data_out = 8'hE7;
                    16'h8BDD: data_out = 8'hE8;
                    16'h8BDE: data_out = 8'hE9;
                    16'h8BDF: data_out = 8'hEA;
                    16'h8BE0: data_out = 8'hEB;
                    16'h8BE1: data_out = 8'hEC;
                    16'h8BE2: data_out = 8'hED;
                    16'h8BE3: data_out = 8'hEE;
                    16'h8BE4: data_out = 8'hEF;
                    16'h8BE5: data_out = 8'hF0;
                    16'h8BE6: data_out = 8'hF1;
                    16'h8BE7: data_out = 8'hF2;
                    16'h8BE8: data_out = 8'hF3;
                    16'h8BE9: data_out = 8'hF4;
                    16'h8BEA: data_out = 8'hF5;
                    16'h8BEB: data_out = 8'hF6;
                    16'h8BEC: data_out = 8'hF7;
                    16'h8BED: data_out = 8'hF8;
                    16'h8BEE: data_out = 8'hF9;
                    16'h8BEF: data_out = 8'hFA;
                    16'h8BF0: data_out = 8'hFB;
                    16'h8BF1: data_out = 8'hFC;
                    16'h8BF2: data_out = 8'hFD;
                    16'h8BF3: data_out = 8'hFE;
                    16'h8BF4: data_out = 8'hFF;
                    16'h8BF5: data_out = 8'h80;
                    16'h8BF6: data_out = 8'h81;
                    16'h8BF7: data_out = 8'h82;
                    16'h8BF8: data_out = 8'h83;
                    16'h8BF9: data_out = 8'h84;
                    16'h8BFA: data_out = 8'h85;
                    16'h8BFB: data_out = 8'h86;
                    16'h8BFC: data_out = 8'h87;
                    16'h8BFD: data_out = 8'h88;
                    16'h8BFE: data_out = 8'h89;
                    16'h8BFF: data_out = 8'h8A;
                    16'h8C00: data_out = 8'h8C;
                    16'h8C01: data_out = 8'h8B;
                    16'h8C02: data_out = 8'h8A;
                    16'h8C03: data_out = 8'h89;
                    16'h8C04: data_out = 8'h88;
                    16'h8C05: data_out = 8'h87;
                    16'h8C06: data_out = 8'h86;
                    16'h8C07: data_out = 8'h85;
                    16'h8C08: data_out = 8'h84;
                    16'h8C09: data_out = 8'h83;
                    16'h8C0A: data_out = 8'h82;
                    16'h8C0B: data_out = 8'h81;
                    16'h8C0C: data_out = 8'h0;
                    16'h8C0D: data_out = 8'h1;
                    16'h8C0E: data_out = 8'h2;
                    16'h8C0F: data_out = 8'h3;
                    16'h8C10: data_out = 8'h4;
                    16'h8C11: data_out = 8'h5;
                    16'h8C12: data_out = 8'h6;
                    16'h8C13: data_out = 8'h7;
                    16'h8C14: data_out = 8'h8;
                    16'h8C15: data_out = 8'h9;
                    16'h8C16: data_out = 8'hA;
                    16'h8C17: data_out = 8'hB;
                    16'h8C18: data_out = 8'hC;
                    16'h8C19: data_out = 8'hD;
                    16'h8C1A: data_out = 8'hE;
                    16'h8C1B: data_out = 8'hF;
                    16'h8C1C: data_out = 8'h10;
                    16'h8C1D: data_out = 8'h11;
                    16'h8C1E: data_out = 8'h12;
                    16'h8C1F: data_out = 8'h13;
                    16'h8C20: data_out = 8'h14;
                    16'h8C21: data_out = 8'h15;
                    16'h8C22: data_out = 8'h16;
                    16'h8C23: data_out = 8'h17;
                    16'h8C24: data_out = 8'h18;
                    16'h8C25: data_out = 8'h19;
                    16'h8C26: data_out = 8'h1A;
                    16'h8C27: data_out = 8'h1B;
                    16'h8C28: data_out = 8'h1C;
                    16'h8C29: data_out = 8'h1D;
                    16'h8C2A: data_out = 8'h1E;
                    16'h8C2B: data_out = 8'h1F;
                    16'h8C2C: data_out = 8'h20;
                    16'h8C2D: data_out = 8'h21;
                    16'h8C2E: data_out = 8'h22;
                    16'h8C2F: data_out = 8'h23;
                    16'h8C30: data_out = 8'h24;
                    16'h8C31: data_out = 8'h25;
                    16'h8C32: data_out = 8'h26;
                    16'h8C33: data_out = 8'h27;
                    16'h8C34: data_out = 8'h28;
                    16'h8C35: data_out = 8'h29;
                    16'h8C36: data_out = 8'h2A;
                    16'h8C37: data_out = 8'h2B;
                    16'h8C38: data_out = 8'h2C;
                    16'h8C39: data_out = 8'h2D;
                    16'h8C3A: data_out = 8'h2E;
                    16'h8C3B: data_out = 8'h2F;
                    16'h8C3C: data_out = 8'h30;
                    16'h8C3D: data_out = 8'h31;
                    16'h8C3E: data_out = 8'h32;
                    16'h8C3F: data_out = 8'h33;
                    16'h8C40: data_out = 8'h34;
                    16'h8C41: data_out = 8'h35;
                    16'h8C42: data_out = 8'h36;
                    16'h8C43: data_out = 8'h37;
                    16'h8C44: data_out = 8'h38;
                    16'h8C45: data_out = 8'h39;
                    16'h8C46: data_out = 8'h3A;
                    16'h8C47: data_out = 8'h3B;
                    16'h8C48: data_out = 8'h3C;
                    16'h8C49: data_out = 8'h3D;
                    16'h8C4A: data_out = 8'h3E;
                    16'h8C4B: data_out = 8'h3F;
                    16'h8C4C: data_out = 8'h40;
                    16'h8C4D: data_out = 8'h41;
                    16'h8C4E: data_out = 8'h42;
                    16'h8C4F: data_out = 8'h43;
                    16'h8C50: data_out = 8'h44;
                    16'h8C51: data_out = 8'h45;
                    16'h8C52: data_out = 8'h46;
                    16'h8C53: data_out = 8'h47;
                    16'h8C54: data_out = 8'h48;
                    16'h8C55: data_out = 8'h49;
                    16'h8C56: data_out = 8'h4A;
                    16'h8C57: data_out = 8'h4B;
                    16'h8C58: data_out = 8'h4C;
                    16'h8C59: data_out = 8'h4D;
                    16'h8C5A: data_out = 8'h4E;
                    16'h8C5B: data_out = 8'h4F;
                    16'h8C5C: data_out = 8'h50;
                    16'h8C5D: data_out = 8'h51;
                    16'h8C5E: data_out = 8'h52;
                    16'h8C5F: data_out = 8'h53;
                    16'h8C60: data_out = 8'h54;
                    16'h8C61: data_out = 8'h55;
                    16'h8C62: data_out = 8'h56;
                    16'h8C63: data_out = 8'h57;
                    16'h8C64: data_out = 8'h58;
                    16'h8C65: data_out = 8'h59;
                    16'h8C66: data_out = 8'h5A;
                    16'h8C67: data_out = 8'h5B;
                    16'h8C68: data_out = 8'h5C;
                    16'h8C69: data_out = 8'h5D;
                    16'h8C6A: data_out = 8'h5E;
                    16'h8C6B: data_out = 8'h5F;
                    16'h8C6C: data_out = 8'h60;
                    16'h8C6D: data_out = 8'h61;
                    16'h8C6E: data_out = 8'h62;
                    16'h8C6F: data_out = 8'h63;
                    16'h8C70: data_out = 8'h64;
                    16'h8C71: data_out = 8'h65;
                    16'h8C72: data_out = 8'h66;
                    16'h8C73: data_out = 8'h67;
                    16'h8C74: data_out = 8'h68;
                    16'h8C75: data_out = 8'h69;
                    16'h8C76: data_out = 8'h6A;
                    16'h8C77: data_out = 8'h6B;
                    16'h8C78: data_out = 8'h6C;
                    16'h8C79: data_out = 8'h6D;
                    16'h8C7A: data_out = 8'h6E;
                    16'h8C7B: data_out = 8'h6F;
                    16'h8C7C: data_out = 8'h70;
                    16'h8C7D: data_out = 8'h71;
                    16'h8C7E: data_out = 8'h72;
                    16'h8C7F: data_out = 8'h73;
                    16'h8C80: data_out = 8'h8C;
                    16'h8C81: data_out = 8'h8D;
                    16'h8C82: data_out = 8'h8E;
                    16'h8C83: data_out = 8'h8F;
                    16'h8C84: data_out = 8'h90;
                    16'h8C85: data_out = 8'h91;
                    16'h8C86: data_out = 8'h92;
                    16'h8C87: data_out = 8'h93;
                    16'h8C88: data_out = 8'h94;
                    16'h8C89: data_out = 8'h95;
                    16'h8C8A: data_out = 8'h96;
                    16'h8C8B: data_out = 8'h97;
                    16'h8C8C: data_out = 8'h98;
                    16'h8C8D: data_out = 8'h99;
                    16'h8C8E: data_out = 8'h9A;
                    16'h8C8F: data_out = 8'h9B;
                    16'h8C90: data_out = 8'h9C;
                    16'h8C91: data_out = 8'h9D;
                    16'h8C92: data_out = 8'h9E;
                    16'h8C93: data_out = 8'h9F;
                    16'h8C94: data_out = 8'hA0;
                    16'h8C95: data_out = 8'hA1;
                    16'h8C96: data_out = 8'hA2;
                    16'h8C97: data_out = 8'hA3;
                    16'h8C98: data_out = 8'hA4;
                    16'h8C99: data_out = 8'hA5;
                    16'h8C9A: data_out = 8'hA6;
                    16'h8C9B: data_out = 8'hA7;
                    16'h8C9C: data_out = 8'hA8;
                    16'h8C9D: data_out = 8'hA9;
                    16'h8C9E: data_out = 8'hAA;
                    16'h8C9F: data_out = 8'hAB;
                    16'h8CA0: data_out = 8'hAC;
                    16'h8CA1: data_out = 8'hAD;
                    16'h8CA2: data_out = 8'hAE;
                    16'h8CA3: data_out = 8'hAF;
                    16'h8CA4: data_out = 8'hB0;
                    16'h8CA5: data_out = 8'hB1;
                    16'h8CA6: data_out = 8'hB2;
                    16'h8CA7: data_out = 8'hB3;
                    16'h8CA8: data_out = 8'hB4;
                    16'h8CA9: data_out = 8'hB5;
                    16'h8CAA: data_out = 8'hB6;
                    16'h8CAB: data_out = 8'hB7;
                    16'h8CAC: data_out = 8'hB8;
                    16'h8CAD: data_out = 8'hB9;
                    16'h8CAE: data_out = 8'hBA;
                    16'h8CAF: data_out = 8'hBB;
                    16'h8CB0: data_out = 8'hBC;
                    16'h8CB1: data_out = 8'hBD;
                    16'h8CB2: data_out = 8'hBE;
                    16'h8CB3: data_out = 8'hBF;
                    16'h8CB4: data_out = 8'hC0;
                    16'h8CB5: data_out = 8'hC1;
                    16'h8CB6: data_out = 8'hC2;
                    16'h8CB7: data_out = 8'hC3;
                    16'h8CB8: data_out = 8'hC4;
                    16'h8CB9: data_out = 8'hC5;
                    16'h8CBA: data_out = 8'hC6;
                    16'h8CBB: data_out = 8'hC7;
                    16'h8CBC: data_out = 8'hC8;
                    16'h8CBD: data_out = 8'hC9;
                    16'h8CBE: data_out = 8'hCA;
                    16'h8CBF: data_out = 8'hCB;
                    16'h8CC0: data_out = 8'hCC;
                    16'h8CC1: data_out = 8'hCD;
                    16'h8CC2: data_out = 8'hCE;
                    16'h8CC3: data_out = 8'hCF;
                    16'h8CC4: data_out = 8'hD0;
                    16'h8CC5: data_out = 8'hD1;
                    16'h8CC6: data_out = 8'hD2;
                    16'h8CC7: data_out = 8'hD3;
                    16'h8CC8: data_out = 8'hD4;
                    16'h8CC9: data_out = 8'hD5;
                    16'h8CCA: data_out = 8'hD6;
                    16'h8CCB: data_out = 8'hD7;
                    16'h8CCC: data_out = 8'hD8;
                    16'h8CCD: data_out = 8'hD9;
                    16'h8CCE: data_out = 8'hDA;
                    16'h8CCF: data_out = 8'hDB;
                    16'h8CD0: data_out = 8'hDC;
                    16'h8CD1: data_out = 8'hDD;
                    16'h8CD2: data_out = 8'hDE;
                    16'h8CD3: data_out = 8'hDF;
                    16'h8CD4: data_out = 8'hE0;
                    16'h8CD5: data_out = 8'hE1;
                    16'h8CD6: data_out = 8'hE2;
                    16'h8CD7: data_out = 8'hE3;
                    16'h8CD8: data_out = 8'hE4;
                    16'h8CD9: data_out = 8'hE5;
                    16'h8CDA: data_out = 8'hE6;
                    16'h8CDB: data_out = 8'hE7;
                    16'h8CDC: data_out = 8'hE8;
                    16'h8CDD: data_out = 8'hE9;
                    16'h8CDE: data_out = 8'hEA;
                    16'h8CDF: data_out = 8'hEB;
                    16'h8CE0: data_out = 8'hEC;
                    16'h8CE1: data_out = 8'hED;
                    16'h8CE2: data_out = 8'hEE;
                    16'h8CE3: data_out = 8'hEF;
                    16'h8CE4: data_out = 8'hF0;
                    16'h8CE5: data_out = 8'hF1;
                    16'h8CE6: data_out = 8'hF2;
                    16'h8CE7: data_out = 8'hF3;
                    16'h8CE8: data_out = 8'hF4;
                    16'h8CE9: data_out = 8'hF5;
                    16'h8CEA: data_out = 8'hF6;
                    16'h8CEB: data_out = 8'hF7;
                    16'h8CEC: data_out = 8'hF8;
                    16'h8CED: data_out = 8'hF9;
                    16'h8CEE: data_out = 8'hFA;
                    16'h8CEF: data_out = 8'hFB;
                    16'h8CF0: data_out = 8'hFC;
                    16'h8CF1: data_out = 8'hFD;
                    16'h8CF2: data_out = 8'hFE;
                    16'h8CF3: data_out = 8'hFF;
                    16'h8CF4: data_out = 8'h80;
                    16'h8CF5: data_out = 8'h81;
                    16'h8CF6: data_out = 8'h82;
                    16'h8CF7: data_out = 8'h83;
                    16'h8CF8: data_out = 8'h84;
                    16'h8CF9: data_out = 8'h85;
                    16'h8CFA: data_out = 8'h86;
                    16'h8CFB: data_out = 8'h87;
                    16'h8CFC: data_out = 8'h88;
                    16'h8CFD: data_out = 8'h89;
                    16'h8CFE: data_out = 8'h8A;
                    16'h8CFF: data_out = 8'h8B;
                    16'h8D00: data_out = 8'h8D;
                    16'h8D01: data_out = 8'h8C;
                    16'h8D02: data_out = 8'h8B;
                    16'h8D03: data_out = 8'h8A;
                    16'h8D04: data_out = 8'h89;
                    16'h8D05: data_out = 8'h88;
                    16'h8D06: data_out = 8'h87;
                    16'h8D07: data_out = 8'h86;
                    16'h8D08: data_out = 8'h85;
                    16'h8D09: data_out = 8'h84;
                    16'h8D0A: data_out = 8'h83;
                    16'h8D0B: data_out = 8'h82;
                    16'h8D0C: data_out = 8'h81;
                    16'h8D0D: data_out = 8'h0;
                    16'h8D0E: data_out = 8'h1;
                    16'h8D0F: data_out = 8'h2;
                    16'h8D10: data_out = 8'h3;
                    16'h8D11: data_out = 8'h4;
                    16'h8D12: data_out = 8'h5;
                    16'h8D13: data_out = 8'h6;
                    16'h8D14: data_out = 8'h7;
                    16'h8D15: data_out = 8'h8;
                    16'h8D16: data_out = 8'h9;
                    16'h8D17: data_out = 8'hA;
                    16'h8D18: data_out = 8'hB;
                    16'h8D19: data_out = 8'hC;
                    16'h8D1A: data_out = 8'hD;
                    16'h8D1B: data_out = 8'hE;
                    16'h8D1C: data_out = 8'hF;
                    16'h8D1D: data_out = 8'h10;
                    16'h8D1E: data_out = 8'h11;
                    16'h8D1F: data_out = 8'h12;
                    16'h8D20: data_out = 8'h13;
                    16'h8D21: data_out = 8'h14;
                    16'h8D22: data_out = 8'h15;
                    16'h8D23: data_out = 8'h16;
                    16'h8D24: data_out = 8'h17;
                    16'h8D25: data_out = 8'h18;
                    16'h8D26: data_out = 8'h19;
                    16'h8D27: data_out = 8'h1A;
                    16'h8D28: data_out = 8'h1B;
                    16'h8D29: data_out = 8'h1C;
                    16'h8D2A: data_out = 8'h1D;
                    16'h8D2B: data_out = 8'h1E;
                    16'h8D2C: data_out = 8'h1F;
                    16'h8D2D: data_out = 8'h20;
                    16'h8D2E: data_out = 8'h21;
                    16'h8D2F: data_out = 8'h22;
                    16'h8D30: data_out = 8'h23;
                    16'h8D31: data_out = 8'h24;
                    16'h8D32: data_out = 8'h25;
                    16'h8D33: data_out = 8'h26;
                    16'h8D34: data_out = 8'h27;
                    16'h8D35: data_out = 8'h28;
                    16'h8D36: data_out = 8'h29;
                    16'h8D37: data_out = 8'h2A;
                    16'h8D38: data_out = 8'h2B;
                    16'h8D39: data_out = 8'h2C;
                    16'h8D3A: data_out = 8'h2D;
                    16'h8D3B: data_out = 8'h2E;
                    16'h8D3C: data_out = 8'h2F;
                    16'h8D3D: data_out = 8'h30;
                    16'h8D3E: data_out = 8'h31;
                    16'h8D3F: data_out = 8'h32;
                    16'h8D40: data_out = 8'h33;
                    16'h8D41: data_out = 8'h34;
                    16'h8D42: data_out = 8'h35;
                    16'h8D43: data_out = 8'h36;
                    16'h8D44: data_out = 8'h37;
                    16'h8D45: data_out = 8'h38;
                    16'h8D46: data_out = 8'h39;
                    16'h8D47: data_out = 8'h3A;
                    16'h8D48: data_out = 8'h3B;
                    16'h8D49: data_out = 8'h3C;
                    16'h8D4A: data_out = 8'h3D;
                    16'h8D4B: data_out = 8'h3E;
                    16'h8D4C: data_out = 8'h3F;
                    16'h8D4D: data_out = 8'h40;
                    16'h8D4E: data_out = 8'h41;
                    16'h8D4F: data_out = 8'h42;
                    16'h8D50: data_out = 8'h43;
                    16'h8D51: data_out = 8'h44;
                    16'h8D52: data_out = 8'h45;
                    16'h8D53: data_out = 8'h46;
                    16'h8D54: data_out = 8'h47;
                    16'h8D55: data_out = 8'h48;
                    16'h8D56: data_out = 8'h49;
                    16'h8D57: data_out = 8'h4A;
                    16'h8D58: data_out = 8'h4B;
                    16'h8D59: data_out = 8'h4C;
                    16'h8D5A: data_out = 8'h4D;
                    16'h8D5B: data_out = 8'h4E;
                    16'h8D5C: data_out = 8'h4F;
                    16'h8D5D: data_out = 8'h50;
                    16'h8D5E: data_out = 8'h51;
                    16'h8D5F: data_out = 8'h52;
                    16'h8D60: data_out = 8'h53;
                    16'h8D61: data_out = 8'h54;
                    16'h8D62: data_out = 8'h55;
                    16'h8D63: data_out = 8'h56;
                    16'h8D64: data_out = 8'h57;
                    16'h8D65: data_out = 8'h58;
                    16'h8D66: data_out = 8'h59;
                    16'h8D67: data_out = 8'h5A;
                    16'h8D68: data_out = 8'h5B;
                    16'h8D69: data_out = 8'h5C;
                    16'h8D6A: data_out = 8'h5D;
                    16'h8D6B: data_out = 8'h5E;
                    16'h8D6C: data_out = 8'h5F;
                    16'h8D6D: data_out = 8'h60;
                    16'h8D6E: data_out = 8'h61;
                    16'h8D6F: data_out = 8'h62;
                    16'h8D70: data_out = 8'h63;
                    16'h8D71: data_out = 8'h64;
                    16'h8D72: data_out = 8'h65;
                    16'h8D73: data_out = 8'h66;
                    16'h8D74: data_out = 8'h67;
                    16'h8D75: data_out = 8'h68;
                    16'h8D76: data_out = 8'h69;
                    16'h8D77: data_out = 8'h6A;
                    16'h8D78: data_out = 8'h6B;
                    16'h8D79: data_out = 8'h6C;
                    16'h8D7A: data_out = 8'h6D;
                    16'h8D7B: data_out = 8'h6E;
                    16'h8D7C: data_out = 8'h6F;
                    16'h8D7D: data_out = 8'h70;
                    16'h8D7E: data_out = 8'h71;
                    16'h8D7F: data_out = 8'h72;
                    16'h8D80: data_out = 8'h8D;
                    16'h8D81: data_out = 8'h8E;
                    16'h8D82: data_out = 8'h8F;
                    16'h8D83: data_out = 8'h90;
                    16'h8D84: data_out = 8'h91;
                    16'h8D85: data_out = 8'h92;
                    16'h8D86: data_out = 8'h93;
                    16'h8D87: data_out = 8'h94;
                    16'h8D88: data_out = 8'h95;
                    16'h8D89: data_out = 8'h96;
                    16'h8D8A: data_out = 8'h97;
                    16'h8D8B: data_out = 8'h98;
                    16'h8D8C: data_out = 8'h99;
                    16'h8D8D: data_out = 8'h9A;
                    16'h8D8E: data_out = 8'h9B;
                    16'h8D8F: data_out = 8'h9C;
                    16'h8D90: data_out = 8'h9D;
                    16'h8D91: data_out = 8'h9E;
                    16'h8D92: data_out = 8'h9F;
                    16'h8D93: data_out = 8'hA0;
                    16'h8D94: data_out = 8'hA1;
                    16'h8D95: data_out = 8'hA2;
                    16'h8D96: data_out = 8'hA3;
                    16'h8D97: data_out = 8'hA4;
                    16'h8D98: data_out = 8'hA5;
                    16'h8D99: data_out = 8'hA6;
                    16'h8D9A: data_out = 8'hA7;
                    16'h8D9B: data_out = 8'hA8;
                    16'h8D9C: data_out = 8'hA9;
                    16'h8D9D: data_out = 8'hAA;
                    16'h8D9E: data_out = 8'hAB;
                    16'h8D9F: data_out = 8'hAC;
                    16'h8DA0: data_out = 8'hAD;
                    16'h8DA1: data_out = 8'hAE;
                    16'h8DA2: data_out = 8'hAF;
                    16'h8DA3: data_out = 8'hB0;
                    16'h8DA4: data_out = 8'hB1;
                    16'h8DA5: data_out = 8'hB2;
                    16'h8DA6: data_out = 8'hB3;
                    16'h8DA7: data_out = 8'hB4;
                    16'h8DA8: data_out = 8'hB5;
                    16'h8DA9: data_out = 8'hB6;
                    16'h8DAA: data_out = 8'hB7;
                    16'h8DAB: data_out = 8'hB8;
                    16'h8DAC: data_out = 8'hB9;
                    16'h8DAD: data_out = 8'hBA;
                    16'h8DAE: data_out = 8'hBB;
                    16'h8DAF: data_out = 8'hBC;
                    16'h8DB0: data_out = 8'hBD;
                    16'h8DB1: data_out = 8'hBE;
                    16'h8DB2: data_out = 8'hBF;
                    16'h8DB3: data_out = 8'hC0;
                    16'h8DB4: data_out = 8'hC1;
                    16'h8DB5: data_out = 8'hC2;
                    16'h8DB6: data_out = 8'hC3;
                    16'h8DB7: data_out = 8'hC4;
                    16'h8DB8: data_out = 8'hC5;
                    16'h8DB9: data_out = 8'hC6;
                    16'h8DBA: data_out = 8'hC7;
                    16'h8DBB: data_out = 8'hC8;
                    16'h8DBC: data_out = 8'hC9;
                    16'h8DBD: data_out = 8'hCA;
                    16'h8DBE: data_out = 8'hCB;
                    16'h8DBF: data_out = 8'hCC;
                    16'h8DC0: data_out = 8'hCD;
                    16'h8DC1: data_out = 8'hCE;
                    16'h8DC2: data_out = 8'hCF;
                    16'h8DC3: data_out = 8'hD0;
                    16'h8DC4: data_out = 8'hD1;
                    16'h8DC5: data_out = 8'hD2;
                    16'h8DC6: data_out = 8'hD3;
                    16'h8DC7: data_out = 8'hD4;
                    16'h8DC8: data_out = 8'hD5;
                    16'h8DC9: data_out = 8'hD6;
                    16'h8DCA: data_out = 8'hD7;
                    16'h8DCB: data_out = 8'hD8;
                    16'h8DCC: data_out = 8'hD9;
                    16'h8DCD: data_out = 8'hDA;
                    16'h8DCE: data_out = 8'hDB;
                    16'h8DCF: data_out = 8'hDC;
                    16'h8DD0: data_out = 8'hDD;
                    16'h8DD1: data_out = 8'hDE;
                    16'h8DD2: data_out = 8'hDF;
                    16'h8DD3: data_out = 8'hE0;
                    16'h8DD4: data_out = 8'hE1;
                    16'h8DD5: data_out = 8'hE2;
                    16'h8DD6: data_out = 8'hE3;
                    16'h8DD7: data_out = 8'hE4;
                    16'h8DD8: data_out = 8'hE5;
                    16'h8DD9: data_out = 8'hE6;
                    16'h8DDA: data_out = 8'hE7;
                    16'h8DDB: data_out = 8'hE8;
                    16'h8DDC: data_out = 8'hE9;
                    16'h8DDD: data_out = 8'hEA;
                    16'h8DDE: data_out = 8'hEB;
                    16'h8DDF: data_out = 8'hEC;
                    16'h8DE0: data_out = 8'hED;
                    16'h8DE1: data_out = 8'hEE;
                    16'h8DE2: data_out = 8'hEF;
                    16'h8DE3: data_out = 8'hF0;
                    16'h8DE4: data_out = 8'hF1;
                    16'h8DE5: data_out = 8'hF2;
                    16'h8DE6: data_out = 8'hF3;
                    16'h8DE7: data_out = 8'hF4;
                    16'h8DE8: data_out = 8'hF5;
                    16'h8DE9: data_out = 8'hF6;
                    16'h8DEA: data_out = 8'hF7;
                    16'h8DEB: data_out = 8'hF8;
                    16'h8DEC: data_out = 8'hF9;
                    16'h8DED: data_out = 8'hFA;
                    16'h8DEE: data_out = 8'hFB;
                    16'h8DEF: data_out = 8'hFC;
                    16'h8DF0: data_out = 8'hFD;
                    16'h8DF1: data_out = 8'hFE;
                    16'h8DF2: data_out = 8'hFF;
                    16'h8DF3: data_out = 8'h80;
                    16'h8DF4: data_out = 8'h81;
                    16'h8DF5: data_out = 8'h82;
                    16'h8DF6: data_out = 8'h83;
                    16'h8DF7: data_out = 8'h84;
                    16'h8DF8: data_out = 8'h85;
                    16'h8DF9: data_out = 8'h86;
                    16'h8DFA: data_out = 8'h87;
                    16'h8DFB: data_out = 8'h88;
                    16'h8DFC: data_out = 8'h89;
                    16'h8DFD: data_out = 8'h8A;
                    16'h8DFE: data_out = 8'h8B;
                    16'h8DFF: data_out = 8'h8C;
                    16'h8E00: data_out = 8'h8E;
                    16'h8E01: data_out = 8'h8D;
                    16'h8E02: data_out = 8'h8C;
                    16'h8E03: data_out = 8'h8B;
                    16'h8E04: data_out = 8'h8A;
                    16'h8E05: data_out = 8'h89;
                    16'h8E06: data_out = 8'h88;
                    16'h8E07: data_out = 8'h87;
                    16'h8E08: data_out = 8'h86;
                    16'h8E09: data_out = 8'h85;
                    16'h8E0A: data_out = 8'h84;
                    16'h8E0B: data_out = 8'h83;
                    16'h8E0C: data_out = 8'h82;
                    16'h8E0D: data_out = 8'h81;
                    16'h8E0E: data_out = 8'h0;
                    16'h8E0F: data_out = 8'h1;
                    16'h8E10: data_out = 8'h2;
                    16'h8E11: data_out = 8'h3;
                    16'h8E12: data_out = 8'h4;
                    16'h8E13: data_out = 8'h5;
                    16'h8E14: data_out = 8'h6;
                    16'h8E15: data_out = 8'h7;
                    16'h8E16: data_out = 8'h8;
                    16'h8E17: data_out = 8'h9;
                    16'h8E18: data_out = 8'hA;
                    16'h8E19: data_out = 8'hB;
                    16'h8E1A: data_out = 8'hC;
                    16'h8E1B: data_out = 8'hD;
                    16'h8E1C: data_out = 8'hE;
                    16'h8E1D: data_out = 8'hF;
                    16'h8E1E: data_out = 8'h10;
                    16'h8E1F: data_out = 8'h11;
                    16'h8E20: data_out = 8'h12;
                    16'h8E21: data_out = 8'h13;
                    16'h8E22: data_out = 8'h14;
                    16'h8E23: data_out = 8'h15;
                    16'h8E24: data_out = 8'h16;
                    16'h8E25: data_out = 8'h17;
                    16'h8E26: data_out = 8'h18;
                    16'h8E27: data_out = 8'h19;
                    16'h8E28: data_out = 8'h1A;
                    16'h8E29: data_out = 8'h1B;
                    16'h8E2A: data_out = 8'h1C;
                    16'h8E2B: data_out = 8'h1D;
                    16'h8E2C: data_out = 8'h1E;
                    16'h8E2D: data_out = 8'h1F;
                    16'h8E2E: data_out = 8'h20;
                    16'h8E2F: data_out = 8'h21;
                    16'h8E30: data_out = 8'h22;
                    16'h8E31: data_out = 8'h23;
                    16'h8E32: data_out = 8'h24;
                    16'h8E33: data_out = 8'h25;
                    16'h8E34: data_out = 8'h26;
                    16'h8E35: data_out = 8'h27;
                    16'h8E36: data_out = 8'h28;
                    16'h8E37: data_out = 8'h29;
                    16'h8E38: data_out = 8'h2A;
                    16'h8E39: data_out = 8'h2B;
                    16'h8E3A: data_out = 8'h2C;
                    16'h8E3B: data_out = 8'h2D;
                    16'h8E3C: data_out = 8'h2E;
                    16'h8E3D: data_out = 8'h2F;
                    16'h8E3E: data_out = 8'h30;
                    16'h8E3F: data_out = 8'h31;
                    16'h8E40: data_out = 8'h32;
                    16'h8E41: data_out = 8'h33;
                    16'h8E42: data_out = 8'h34;
                    16'h8E43: data_out = 8'h35;
                    16'h8E44: data_out = 8'h36;
                    16'h8E45: data_out = 8'h37;
                    16'h8E46: data_out = 8'h38;
                    16'h8E47: data_out = 8'h39;
                    16'h8E48: data_out = 8'h3A;
                    16'h8E49: data_out = 8'h3B;
                    16'h8E4A: data_out = 8'h3C;
                    16'h8E4B: data_out = 8'h3D;
                    16'h8E4C: data_out = 8'h3E;
                    16'h8E4D: data_out = 8'h3F;
                    16'h8E4E: data_out = 8'h40;
                    16'h8E4F: data_out = 8'h41;
                    16'h8E50: data_out = 8'h42;
                    16'h8E51: data_out = 8'h43;
                    16'h8E52: data_out = 8'h44;
                    16'h8E53: data_out = 8'h45;
                    16'h8E54: data_out = 8'h46;
                    16'h8E55: data_out = 8'h47;
                    16'h8E56: data_out = 8'h48;
                    16'h8E57: data_out = 8'h49;
                    16'h8E58: data_out = 8'h4A;
                    16'h8E59: data_out = 8'h4B;
                    16'h8E5A: data_out = 8'h4C;
                    16'h8E5B: data_out = 8'h4D;
                    16'h8E5C: data_out = 8'h4E;
                    16'h8E5D: data_out = 8'h4F;
                    16'h8E5E: data_out = 8'h50;
                    16'h8E5F: data_out = 8'h51;
                    16'h8E60: data_out = 8'h52;
                    16'h8E61: data_out = 8'h53;
                    16'h8E62: data_out = 8'h54;
                    16'h8E63: data_out = 8'h55;
                    16'h8E64: data_out = 8'h56;
                    16'h8E65: data_out = 8'h57;
                    16'h8E66: data_out = 8'h58;
                    16'h8E67: data_out = 8'h59;
                    16'h8E68: data_out = 8'h5A;
                    16'h8E69: data_out = 8'h5B;
                    16'h8E6A: data_out = 8'h5C;
                    16'h8E6B: data_out = 8'h5D;
                    16'h8E6C: data_out = 8'h5E;
                    16'h8E6D: data_out = 8'h5F;
                    16'h8E6E: data_out = 8'h60;
                    16'h8E6F: data_out = 8'h61;
                    16'h8E70: data_out = 8'h62;
                    16'h8E71: data_out = 8'h63;
                    16'h8E72: data_out = 8'h64;
                    16'h8E73: data_out = 8'h65;
                    16'h8E74: data_out = 8'h66;
                    16'h8E75: data_out = 8'h67;
                    16'h8E76: data_out = 8'h68;
                    16'h8E77: data_out = 8'h69;
                    16'h8E78: data_out = 8'h6A;
                    16'h8E79: data_out = 8'h6B;
                    16'h8E7A: data_out = 8'h6C;
                    16'h8E7B: data_out = 8'h6D;
                    16'h8E7C: data_out = 8'h6E;
                    16'h8E7D: data_out = 8'h6F;
                    16'h8E7E: data_out = 8'h70;
                    16'h8E7F: data_out = 8'h71;
                    16'h8E80: data_out = 8'h8E;
                    16'h8E81: data_out = 8'h8F;
                    16'h8E82: data_out = 8'h90;
                    16'h8E83: data_out = 8'h91;
                    16'h8E84: data_out = 8'h92;
                    16'h8E85: data_out = 8'h93;
                    16'h8E86: data_out = 8'h94;
                    16'h8E87: data_out = 8'h95;
                    16'h8E88: data_out = 8'h96;
                    16'h8E89: data_out = 8'h97;
                    16'h8E8A: data_out = 8'h98;
                    16'h8E8B: data_out = 8'h99;
                    16'h8E8C: data_out = 8'h9A;
                    16'h8E8D: data_out = 8'h9B;
                    16'h8E8E: data_out = 8'h9C;
                    16'h8E8F: data_out = 8'h9D;
                    16'h8E90: data_out = 8'h9E;
                    16'h8E91: data_out = 8'h9F;
                    16'h8E92: data_out = 8'hA0;
                    16'h8E93: data_out = 8'hA1;
                    16'h8E94: data_out = 8'hA2;
                    16'h8E95: data_out = 8'hA3;
                    16'h8E96: data_out = 8'hA4;
                    16'h8E97: data_out = 8'hA5;
                    16'h8E98: data_out = 8'hA6;
                    16'h8E99: data_out = 8'hA7;
                    16'h8E9A: data_out = 8'hA8;
                    16'h8E9B: data_out = 8'hA9;
                    16'h8E9C: data_out = 8'hAA;
                    16'h8E9D: data_out = 8'hAB;
                    16'h8E9E: data_out = 8'hAC;
                    16'h8E9F: data_out = 8'hAD;
                    16'h8EA0: data_out = 8'hAE;
                    16'h8EA1: data_out = 8'hAF;
                    16'h8EA2: data_out = 8'hB0;
                    16'h8EA3: data_out = 8'hB1;
                    16'h8EA4: data_out = 8'hB2;
                    16'h8EA5: data_out = 8'hB3;
                    16'h8EA6: data_out = 8'hB4;
                    16'h8EA7: data_out = 8'hB5;
                    16'h8EA8: data_out = 8'hB6;
                    16'h8EA9: data_out = 8'hB7;
                    16'h8EAA: data_out = 8'hB8;
                    16'h8EAB: data_out = 8'hB9;
                    16'h8EAC: data_out = 8'hBA;
                    16'h8EAD: data_out = 8'hBB;
                    16'h8EAE: data_out = 8'hBC;
                    16'h8EAF: data_out = 8'hBD;
                    16'h8EB0: data_out = 8'hBE;
                    16'h8EB1: data_out = 8'hBF;
                    16'h8EB2: data_out = 8'hC0;
                    16'h8EB3: data_out = 8'hC1;
                    16'h8EB4: data_out = 8'hC2;
                    16'h8EB5: data_out = 8'hC3;
                    16'h8EB6: data_out = 8'hC4;
                    16'h8EB7: data_out = 8'hC5;
                    16'h8EB8: data_out = 8'hC6;
                    16'h8EB9: data_out = 8'hC7;
                    16'h8EBA: data_out = 8'hC8;
                    16'h8EBB: data_out = 8'hC9;
                    16'h8EBC: data_out = 8'hCA;
                    16'h8EBD: data_out = 8'hCB;
                    16'h8EBE: data_out = 8'hCC;
                    16'h8EBF: data_out = 8'hCD;
                    16'h8EC0: data_out = 8'hCE;
                    16'h8EC1: data_out = 8'hCF;
                    16'h8EC2: data_out = 8'hD0;
                    16'h8EC3: data_out = 8'hD1;
                    16'h8EC4: data_out = 8'hD2;
                    16'h8EC5: data_out = 8'hD3;
                    16'h8EC6: data_out = 8'hD4;
                    16'h8EC7: data_out = 8'hD5;
                    16'h8EC8: data_out = 8'hD6;
                    16'h8EC9: data_out = 8'hD7;
                    16'h8ECA: data_out = 8'hD8;
                    16'h8ECB: data_out = 8'hD9;
                    16'h8ECC: data_out = 8'hDA;
                    16'h8ECD: data_out = 8'hDB;
                    16'h8ECE: data_out = 8'hDC;
                    16'h8ECF: data_out = 8'hDD;
                    16'h8ED0: data_out = 8'hDE;
                    16'h8ED1: data_out = 8'hDF;
                    16'h8ED2: data_out = 8'hE0;
                    16'h8ED3: data_out = 8'hE1;
                    16'h8ED4: data_out = 8'hE2;
                    16'h8ED5: data_out = 8'hE3;
                    16'h8ED6: data_out = 8'hE4;
                    16'h8ED7: data_out = 8'hE5;
                    16'h8ED8: data_out = 8'hE6;
                    16'h8ED9: data_out = 8'hE7;
                    16'h8EDA: data_out = 8'hE8;
                    16'h8EDB: data_out = 8'hE9;
                    16'h8EDC: data_out = 8'hEA;
                    16'h8EDD: data_out = 8'hEB;
                    16'h8EDE: data_out = 8'hEC;
                    16'h8EDF: data_out = 8'hED;
                    16'h8EE0: data_out = 8'hEE;
                    16'h8EE1: data_out = 8'hEF;
                    16'h8EE2: data_out = 8'hF0;
                    16'h8EE3: data_out = 8'hF1;
                    16'h8EE4: data_out = 8'hF2;
                    16'h8EE5: data_out = 8'hF3;
                    16'h8EE6: data_out = 8'hF4;
                    16'h8EE7: data_out = 8'hF5;
                    16'h8EE8: data_out = 8'hF6;
                    16'h8EE9: data_out = 8'hF7;
                    16'h8EEA: data_out = 8'hF8;
                    16'h8EEB: data_out = 8'hF9;
                    16'h8EEC: data_out = 8'hFA;
                    16'h8EED: data_out = 8'hFB;
                    16'h8EEE: data_out = 8'hFC;
                    16'h8EEF: data_out = 8'hFD;
                    16'h8EF0: data_out = 8'hFE;
                    16'h8EF1: data_out = 8'hFF;
                    16'h8EF2: data_out = 8'h80;
                    16'h8EF3: data_out = 8'h81;
                    16'h8EF4: data_out = 8'h82;
                    16'h8EF5: data_out = 8'h83;
                    16'h8EF6: data_out = 8'h84;
                    16'h8EF7: data_out = 8'h85;
                    16'h8EF8: data_out = 8'h86;
                    16'h8EF9: data_out = 8'h87;
                    16'h8EFA: data_out = 8'h88;
                    16'h8EFB: data_out = 8'h89;
                    16'h8EFC: data_out = 8'h8A;
                    16'h8EFD: data_out = 8'h8B;
                    16'h8EFE: data_out = 8'h8C;
                    16'h8EFF: data_out = 8'h8D;
                    16'h8F00: data_out = 8'h8F;
                    16'h8F01: data_out = 8'h8E;
                    16'h8F02: data_out = 8'h8D;
                    16'h8F03: data_out = 8'h8C;
                    16'h8F04: data_out = 8'h8B;
                    16'h8F05: data_out = 8'h8A;
                    16'h8F06: data_out = 8'h89;
                    16'h8F07: data_out = 8'h88;
                    16'h8F08: data_out = 8'h87;
                    16'h8F09: data_out = 8'h86;
                    16'h8F0A: data_out = 8'h85;
                    16'h8F0B: data_out = 8'h84;
                    16'h8F0C: data_out = 8'h83;
                    16'h8F0D: data_out = 8'h82;
                    16'h8F0E: data_out = 8'h81;
                    16'h8F0F: data_out = 8'h0;
                    16'h8F10: data_out = 8'h1;
                    16'h8F11: data_out = 8'h2;
                    16'h8F12: data_out = 8'h3;
                    16'h8F13: data_out = 8'h4;
                    16'h8F14: data_out = 8'h5;
                    16'h8F15: data_out = 8'h6;
                    16'h8F16: data_out = 8'h7;
                    16'h8F17: data_out = 8'h8;
                    16'h8F18: data_out = 8'h9;
                    16'h8F19: data_out = 8'hA;
                    16'h8F1A: data_out = 8'hB;
                    16'h8F1B: data_out = 8'hC;
                    16'h8F1C: data_out = 8'hD;
                    16'h8F1D: data_out = 8'hE;
                    16'h8F1E: data_out = 8'hF;
                    16'h8F1F: data_out = 8'h10;
                    16'h8F20: data_out = 8'h11;
                    16'h8F21: data_out = 8'h12;
                    16'h8F22: data_out = 8'h13;
                    16'h8F23: data_out = 8'h14;
                    16'h8F24: data_out = 8'h15;
                    16'h8F25: data_out = 8'h16;
                    16'h8F26: data_out = 8'h17;
                    16'h8F27: data_out = 8'h18;
                    16'h8F28: data_out = 8'h19;
                    16'h8F29: data_out = 8'h1A;
                    16'h8F2A: data_out = 8'h1B;
                    16'h8F2B: data_out = 8'h1C;
                    16'h8F2C: data_out = 8'h1D;
                    16'h8F2D: data_out = 8'h1E;
                    16'h8F2E: data_out = 8'h1F;
                    16'h8F2F: data_out = 8'h20;
                    16'h8F30: data_out = 8'h21;
                    16'h8F31: data_out = 8'h22;
                    16'h8F32: data_out = 8'h23;
                    16'h8F33: data_out = 8'h24;
                    16'h8F34: data_out = 8'h25;
                    16'h8F35: data_out = 8'h26;
                    16'h8F36: data_out = 8'h27;
                    16'h8F37: data_out = 8'h28;
                    16'h8F38: data_out = 8'h29;
                    16'h8F39: data_out = 8'h2A;
                    16'h8F3A: data_out = 8'h2B;
                    16'h8F3B: data_out = 8'h2C;
                    16'h8F3C: data_out = 8'h2D;
                    16'h8F3D: data_out = 8'h2E;
                    16'h8F3E: data_out = 8'h2F;
                    16'h8F3F: data_out = 8'h30;
                    16'h8F40: data_out = 8'h31;
                    16'h8F41: data_out = 8'h32;
                    16'h8F42: data_out = 8'h33;
                    16'h8F43: data_out = 8'h34;
                    16'h8F44: data_out = 8'h35;
                    16'h8F45: data_out = 8'h36;
                    16'h8F46: data_out = 8'h37;
                    16'h8F47: data_out = 8'h38;
                    16'h8F48: data_out = 8'h39;
                    16'h8F49: data_out = 8'h3A;
                    16'h8F4A: data_out = 8'h3B;
                    16'h8F4B: data_out = 8'h3C;
                    16'h8F4C: data_out = 8'h3D;
                    16'h8F4D: data_out = 8'h3E;
                    16'h8F4E: data_out = 8'h3F;
                    16'h8F4F: data_out = 8'h40;
                    16'h8F50: data_out = 8'h41;
                    16'h8F51: data_out = 8'h42;
                    16'h8F52: data_out = 8'h43;
                    16'h8F53: data_out = 8'h44;
                    16'h8F54: data_out = 8'h45;
                    16'h8F55: data_out = 8'h46;
                    16'h8F56: data_out = 8'h47;
                    16'h8F57: data_out = 8'h48;
                    16'h8F58: data_out = 8'h49;
                    16'h8F59: data_out = 8'h4A;
                    16'h8F5A: data_out = 8'h4B;
                    16'h8F5B: data_out = 8'h4C;
                    16'h8F5C: data_out = 8'h4D;
                    16'h8F5D: data_out = 8'h4E;
                    16'h8F5E: data_out = 8'h4F;
                    16'h8F5F: data_out = 8'h50;
                    16'h8F60: data_out = 8'h51;
                    16'h8F61: data_out = 8'h52;
                    16'h8F62: data_out = 8'h53;
                    16'h8F63: data_out = 8'h54;
                    16'h8F64: data_out = 8'h55;
                    16'h8F65: data_out = 8'h56;
                    16'h8F66: data_out = 8'h57;
                    16'h8F67: data_out = 8'h58;
                    16'h8F68: data_out = 8'h59;
                    16'h8F69: data_out = 8'h5A;
                    16'h8F6A: data_out = 8'h5B;
                    16'h8F6B: data_out = 8'h5C;
                    16'h8F6C: data_out = 8'h5D;
                    16'h8F6D: data_out = 8'h5E;
                    16'h8F6E: data_out = 8'h5F;
                    16'h8F6F: data_out = 8'h60;
                    16'h8F70: data_out = 8'h61;
                    16'h8F71: data_out = 8'h62;
                    16'h8F72: data_out = 8'h63;
                    16'h8F73: data_out = 8'h64;
                    16'h8F74: data_out = 8'h65;
                    16'h8F75: data_out = 8'h66;
                    16'h8F76: data_out = 8'h67;
                    16'h8F77: data_out = 8'h68;
                    16'h8F78: data_out = 8'h69;
                    16'h8F79: data_out = 8'h6A;
                    16'h8F7A: data_out = 8'h6B;
                    16'h8F7B: data_out = 8'h6C;
                    16'h8F7C: data_out = 8'h6D;
                    16'h8F7D: data_out = 8'h6E;
                    16'h8F7E: data_out = 8'h6F;
                    16'h8F7F: data_out = 8'h70;
                    16'h8F80: data_out = 8'h8F;
                    16'h8F81: data_out = 8'h90;
                    16'h8F82: data_out = 8'h91;
                    16'h8F83: data_out = 8'h92;
                    16'h8F84: data_out = 8'h93;
                    16'h8F85: data_out = 8'h94;
                    16'h8F86: data_out = 8'h95;
                    16'h8F87: data_out = 8'h96;
                    16'h8F88: data_out = 8'h97;
                    16'h8F89: data_out = 8'h98;
                    16'h8F8A: data_out = 8'h99;
                    16'h8F8B: data_out = 8'h9A;
                    16'h8F8C: data_out = 8'h9B;
                    16'h8F8D: data_out = 8'h9C;
                    16'h8F8E: data_out = 8'h9D;
                    16'h8F8F: data_out = 8'h9E;
                    16'h8F90: data_out = 8'h9F;
                    16'h8F91: data_out = 8'hA0;
                    16'h8F92: data_out = 8'hA1;
                    16'h8F93: data_out = 8'hA2;
                    16'h8F94: data_out = 8'hA3;
                    16'h8F95: data_out = 8'hA4;
                    16'h8F96: data_out = 8'hA5;
                    16'h8F97: data_out = 8'hA6;
                    16'h8F98: data_out = 8'hA7;
                    16'h8F99: data_out = 8'hA8;
                    16'h8F9A: data_out = 8'hA9;
                    16'h8F9B: data_out = 8'hAA;
                    16'h8F9C: data_out = 8'hAB;
                    16'h8F9D: data_out = 8'hAC;
                    16'h8F9E: data_out = 8'hAD;
                    16'h8F9F: data_out = 8'hAE;
                    16'h8FA0: data_out = 8'hAF;
                    16'h8FA1: data_out = 8'hB0;
                    16'h8FA2: data_out = 8'hB1;
                    16'h8FA3: data_out = 8'hB2;
                    16'h8FA4: data_out = 8'hB3;
                    16'h8FA5: data_out = 8'hB4;
                    16'h8FA6: data_out = 8'hB5;
                    16'h8FA7: data_out = 8'hB6;
                    16'h8FA8: data_out = 8'hB7;
                    16'h8FA9: data_out = 8'hB8;
                    16'h8FAA: data_out = 8'hB9;
                    16'h8FAB: data_out = 8'hBA;
                    16'h8FAC: data_out = 8'hBB;
                    16'h8FAD: data_out = 8'hBC;
                    16'h8FAE: data_out = 8'hBD;
                    16'h8FAF: data_out = 8'hBE;
                    16'h8FB0: data_out = 8'hBF;
                    16'h8FB1: data_out = 8'hC0;
                    16'h8FB2: data_out = 8'hC1;
                    16'h8FB3: data_out = 8'hC2;
                    16'h8FB4: data_out = 8'hC3;
                    16'h8FB5: data_out = 8'hC4;
                    16'h8FB6: data_out = 8'hC5;
                    16'h8FB7: data_out = 8'hC6;
                    16'h8FB8: data_out = 8'hC7;
                    16'h8FB9: data_out = 8'hC8;
                    16'h8FBA: data_out = 8'hC9;
                    16'h8FBB: data_out = 8'hCA;
                    16'h8FBC: data_out = 8'hCB;
                    16'h8FBD: data_out = 8'hCC;
                    16'h8FBE: data_out = 8'hCD;
                    16'h8FBF: data_out = 8'hCE;
                    16'h8FC0: data_out = 8'hCF;
                    16'h8FC1: data_out = 8'hD0;
                    16'h8FC2: data_out = 8'hD1;
                    16'h8FC3: data_out = 8'hD2;
                    16'h8FC4: data_out = 8'hD3;
                    16'h8FC5: data_out = 8'hD4;
                    16'h8FC6: data_out = 8'hD5;
                    16'h8FC7: data_out = 8'hD6;
                    16'h8FC8: data_out = 8'hD7;
                    16'h8FC9: data_out = 8'hD8;
                    16'h8FCA: data_out = 8'hD9;
                    16'h8FCB: data_out = 8'hDA;
                    16'h8FCC: data_out = 8'hDB;
                    16'h8FCD: data_out = 8'hDC;
                    16'h8FCE: data_out = 8'hDD;
                    16'h8FCF: data_out = 8'hDE;
                    16'h8FD0: data_out = 8'hDF;
                    16'h8FD1: data_out = 8'hE0;
                    16'h8FD2: data_out = 8'hE1;
                    16'h8FD3: data_out = 8'hE2;
                    16'h8FD4: data_out = 8'hE3;
                    16'h8FD5: data_out = 8'hE4;
                    16'h8FD6: data_out = 8'hE5;
                    16'h8FD7: data_out = 8'hE6;
                    16'h8FD8: data_out = 8'hE7;
                    16'h8FD9: data_out = 8'hE8;
                    16'h8FDA: data_out = 8'hE9;
                    16'h8FDB: data_out = 8'hEA;
                    16'h8FDC: data_out = 8'hEB;
                    16'h8FDD: data_out = 8'hEC;
                    16'h8FDE: data_out = 8'hED;
                    16'h8FDF: data_out = 8'hEE;
                    16'h8FE0: data_out = 8'hEF;
                    16'h8FE1: data_out = 8'hF0;
                    16'h8FE2: data_out = 8'hF1;
                    16'h8FE3: data_out = 8'hF2;
                    16'h8FE4: data_out = 8'hF3;
                    16'h8FE5: data_out = 8'hF4;
                    16'h8FE6: data_out = 8'hF5;
                    16'h8FE7: data_out = 8'hF6;
                    16'h8FE8: data_out = 8'hF7;
                    16'h8FE9: data_out = 8'hF8;
                    16'h8FEA: data_out = 8'hF9;
                    16'h8FEB: data_out = 8'hFA;
                    16'h8FEC: data_out = 8'hFB;
                    16'h8FED: data_out = 8'hFC;
                    16'h8FEE: data_out = 8'hFD;
                    16'h8FEF: data_out = 8'hFE;
                    16'h8FF0: data_out = 8'hFF;
                    16'h8FF1: data_out = 8'h80;
                    16'h8FF2: data_out = 8'h81;
                    16'h8FF3: data_out = 8'h82;
                    16'h8FF4: data_out = 8'h83;
                    16'h8FF5: data_out = 8'h84;
                    16'h8FF6: data_out = 8'h85;
                    16'h8FF7: data_out = 8'h86;
                    16'h8FF8: data_out = 8'h87;
                    16'h8FF9: data_out = 8'h88;
                    16'h8FFA: data_out = 8'h89;
                    16'h8FFB: data_out = 8'h8A;
                    16'h8FFC: data_out = 8'h8B;
                    16'h8FFD: data_out = 8'h8C;
                    16'h8FFE: data_out = 8'h8D;
                    16'h8FFF: data_out = 8'h8E;
                    16'h9000: data_out = 8'h90;
                    16'h9001: data_out = 8'h8F;
                    16'h9002: data_out = 8'h8E;
                    16'h9003: data_out = 8'h8D;
                    16'h9004: data_out = 8'h8C;
                    16'h9005: data_out = 8'h8B;
                    16'h9006: data_out = 8'h8A;
                    16'h9007: data_out = 8'h89;
                    16'h9008: data_out = 8'h88;
                    16'h9009: data_out = 8'h87;
                    16'h900A: data_out = 8'h86;
                    16'h900B: data_out = 8'h85;
                    16'h900C: data_out = 8'h84;
                    16'h900D: data_out = 8'h83;
                    16'h900E: data_out = 8'h82;
                    16'h900F: data_out = 8'h81;
                    16'h9010: data_out = 8'h0;
                    16'h9011: data_out = 8'h1;
                    16'h9012: data_out = 8'h2;
                    16'h9013: data_out = 8'h3;
                    16'h9014: data_out = 8'h4;
                    16'h9015: data_out = 8'h5;
                    16'h9016: data_out = 8'h6;
                    16'h9017: data_out = 8'h7;
                    16'h9018: data_out = 8'h8;
                    16'h9019: data_out = 8'h9;
                    16'h901A: data_out = 8'hA;
                    16'h901B: data_out = 8'hB;
                    16'h901C: data_out = 8'hC;
                    16'h901D: data_out = 8'hD;
                    16'h901E: data_out = 8'hE;
                    16'h901F: data_out = 8'hF;
                    16'h9020: data_out = 8'h10;
                    16'h9021: data_out = 8'h11;
                    16'h9022: data_out = 8'h12;
                    16'h9023: data_out = 8'h13;
                    16'h9024: data_out = 8'h14;
                    16'h9025: data_out = 8'h15;
                    16'h9026: data_out = 8'h16;
                    16'h9027: data_out = 8'h17;
                    16'h9028: data_out = 8'h18;
                    16'h9029: data_out = 8'h19;
                    16'h902A: data_out = 8'h1A;
                    16'h902B: data_out = 8'h1B;
                    16'h902C: data_out = 8'h1C;
                    16'h902D: data_out = 8'h1D;
                    16'h902E: data_out = 8'h1E;
                    16'h902F: data_out = 8'h1F;
                    16'h9030: data_out = 8'h20;
                    16'h9031: data_out = 8'h21;
                    16'h9032: data_out = 8'h22;
                    16'h9033: data_out = 8'h23;
                    16'h9034: data_out = 8'h24;
                    16'h9035: data_out = 8'h25;
                    16'h9036: data_out = 8'h26;
                    16'h9037: data_out = 8'h27;
                    16'h9038: data_out = 8'h28;
                    16'h9039: data_out = 8'h29;
                    16'h903A: data_out = 8'h2A;
                    16'h903B: data_out = 8'h2B;
                    16'h903C: data_out = 8'h2C;
                    16'h903D: data_out = 8'h2D;
                    16'h903E: data_out = 8'h2E;
                    16'h903F: data_out = 8'h2F;
                    16'h9040: data_out = 8'h30;
                    16'h9041: data_out = 8'h31;
                    16'h9042: data_out = 8'h32;
                    16'h9043: data_out = 8'h33;
                    16'h9044: data_out = 8'h34;
                    16'h9045: data_out = 8'h35;
                    16'h9046: data_out = 8'h36;
                    16'h9047: data_out = 8'h37;
                    16'h9048: data_out = 8'h38;
                    16'h9049: data_out = 8'h39;
                    16'h904A: data_out = 8'h3A;
                    16'h904B: data_out = 8'h3B;
                    16'h904C: data_out = 8'h3C;
                    16'h904D: data_out = 8'h3D;
                    16'h904E: data_out = 8'h3E;
                    16'h904F: data_out = 8'h3F;
                    16'h9050: data_out = 8'h40;
                    16'h9051: data_out = 8'h41;
                    16'h9052: data_out = 8'h42;
                    16'h9053: data_out = 8'h43;
                    16'h9054: data_out = 8'h44;
                    16'h9055: data_out = 8'h45;
                    16'h9056: data_out = 8'h46;
                    16'h9057: data_out = 8'h47;
                    16'h9058: data_out = 8'h48;
                    16'h9059: data_out = 8'h49;
                    16'h905A: data_out = 8'h4A;
                    16'h905B: data_out = 8'h4B;
                    16'h905C: data_out = 8'h4C;
                    16'h905D: data_out = 8'h4D;
                    16'h905E: data_out = 8'h4E;
                    16'h905F: data_out = 8'h4F;
                    16'h9060: data_out = 8'h50;
                    16'h9061: data_out = 8'h51;
                    16'h9062: data_out = 8'h52;
                    16'h9063: data_out = 8'h53;
                    16'h9064: data_out = 8'h54;
                    16'h9065: data_out = 8'h55;
                    16'h9066: data_out = 8'h56;
                    16'h9067: data_out = 8'h57;
                    16'h9068: data_out = 8'h58;
                    16'h9069: data_out = 8'h59;
                    16'h906A: data_out = 8'h5A;
                    16'h906B: data_out = 8'h5B;
                    16'h906C: data_out = 8'h5C;
                    16'h906D: data_out = 8'h5D;
                    16'h906E: data_out = 8'h5E;
                    16'h906F: data_out = 8'h5F;
                    16'h9070: data_out = 8'h60;
                    16'h9071: data_out = 8'h61;
                    16'h9072: data_out = 8'h62;
                    16'h9073: data_out = 8'h63;
                    16'h9074: data_out = 8'h64;
                    16'h9075: data_out = 8'h65;
                    16'h9076: data_out = 8'h66;
                    16'h9077: data_out = 8'h67;
                    16'h9078: data_out = 8'h68;
                    16'h9079: data_out = 8'h69;
                    16'h907A: data_out = 8'h6A;
                    16'h907B: data_out = 8'h6B;
                    16'h907C: data_out = 8'h6C;
                    16'h907D: data_out = 8'h6D;
                    16'h907E: data_out = 8'h6E;
                    16'h907F: data_out = 8'h6F;
                    16'h9080: data_out = 8'h90;
                    16'h9081: data_out = 8'h91;
                    16'h9082: data_out = 8'h92;
                    16'h9083: data_out = 8'h93;
                    16'h9084: data_out = 8'h94;
                    16'h9085: data_out = 8'h95;
                    16'h9086: data_out = 8'h96;
                    16'h9087: data_out = 8'h97;
                    16'h9088: data_out = 8'h98;
                    16'h9089: data_out = 8'h99;
                    16'h908A: data_out = 8'h9A;
                    16'h908B: data_out = 8'h9B;
                    16'h908C: data_out = 8'h9C;
                    16'h908D: data_out = 8'h9D;
                    16'h908E: data_out = 8'h9E;
                    16'h908F: data_out = 8'h9F;
                    16'h9090: data_out = 8'hA0;
                    16'h9091: data_out = 8'hA1;
                    16'h9092: data_out = 8'hA2;
                    16'h9093: data_out = 8'hA3;
                    16'h9094: data_out = 8'hA4;
                    16'h9095: data_out = 8'hA5;
                    16'h9096: data_out = 8'hA6;
                    16'h9097: data_out = 8'hA7;
                    16'h9098: data_out = 8'hA8;
                    16'h9099: data_out = 8'hA9;
                    16'h909A: data_out = 8'hAA;
                    16'h909B: data_out = 8'hAB;
                    16'h909C: data_out = 8'hAC;
                    16'h909D: data_out = 8'hAD;
                    16'h909E: data_out = 8'hAE;
                    16'h909F: data_out = 8'hAF;
                    16'h90A0: data_out = 8'hB0;
                    16'h90A1: data_out = 8'hB1;
                    16'h90A2: data_out = 8'hB2;
                    16'h90A3: data_out = 8'hB3;
                    16'h90A4: data_out = 8'hB4;
                    16'h90A5: data_out = 8'hB5;
                    16'h90A6: data_out = 8'hB6;
                    16'h90A7: data_out = 8'hB7;
                    16'h90A8: data_out = 8'hB8;
                    16'h90A9: data_out = 8'hB9;
                    16'h90AA: data_out = 8'hBA;
                    16'h90AB: data_out = 8'hBB;
                    16'h90AC: data_out = 8'hBC;
                    16'h90AD: data_out = 8'hBD;
                    16'h90AE: data_out = 8'hBE;
                    16'h90AF: data_out = 8'hBF;
                    16'h90B0: data_out = 8'hC0;
                    16'h90B1: data_out = 8'hC1;
                    16'h90B2: data_out = 8'hC2;
                    16'h90B3: data_out = 8'hC3;
                    16'h90B4: data_out = 8'hC4;
                    16'h90B5: data_out = 8'hC5;
                    16'h90B6: data_out = 8'hC6;
                    16'h90B7: data_out = 8'hC7;
                    16'h90B8: data_out = 8'hC8;
                    16'h90B9: data_out = 8'hC9;
                    16'h90BA: data_out = 8'hCA;
                    16'h90BB: data_out = 8'hCB;
                    16'h90BC: data_out = 8'hCC;
                    16'h90BD: data_out = 8'hCD;
                    16'h90BE: data_out = 8'hCE;
                    16'h90BF: data_out = 8'hCF;
                    16'h90C0: data_out = 8'hD0;
                    16'h90C1: data_out = 8'hD1;
                    16'h90C2: data_out = 8'hD2;
                    16'h90C3: data_out = 8'hD3;
                    16'h90C4: data_out = 8'hD4;
                    16'h90C5: data_out = 8'hD5;
                    16'h90C6: data_out = 8'hD6;
                    16'h90C7: data_out = 8'hD7;
                    16'h90C8: data_out = 8'hD8;
                    16'h90C9: data_out = 8'hD9;
                    16'h90CA: data_out = 8'hDA;
                    16'h90CB: data_out = 8'hDB;
                    16'h90CC: data_out = 8'hDC;
                    16'h90CD: data_out = 8'hDD;
                    16'h90CE: data_out = 8'hDE;
                    16'h90CF: data_out = 8'hDF;
                    16'h90D0: data_out = 8'hE0;
                    16'h90D1: data_out = 8'hE1;
                    16'h90D2: data_out = 8'hE2;
                    16'h90D3: data_out = 8'hE3;
                    16'h90D4: data_out = 8'hE4;
                    16'h90D5: data_out = 8'hE5;
                    16'h90D6: data_out = 8'hE6;
                    16'h90D7: data_out = 8'hE7;
                    16'h90D8: data_out = 8'hE8;
                    16'h90D9: data_out = 8'hE9;
                    16'h90DA: data_out = 8'hEA;
                    16'h90DB: data_out = 8'hEB;
                    16'h90DC: data_out = 8'hEC;
                    16'h90DD: data_out = 8'hED;
                    16'h90DE: data_out = 8'hEE;
                    16'h90DF: data_out = 8'hEF;
                    16'h90E0: data_out = 8'hF0;
                    16'h90E1: data_out = 8'hF1;
                    16'h90E2: data_out = 8'hF2;
                    16'h90E3: data_out = 8'hF3;
                    16'h90E4: data_out = 8'hF4;
                    16'h90E5: data_out = 8'hF5;
                    16'h90E6: data_out = 8'hF6;
                    16'h90E7: data_out = 8'hF7;
                    16'h90E8: data_out = 8'hF8;
                    16'h90E9: data_out = 8'hF9;
                    16'h90EA: data_out = 8'hFA;
                    16'h90EB: data_out = 8'hFB;
                    16'h90EC: data_out = 8'hFC;
                    16'h90ED: data_out = 8'hFD;
                    16'h90EE: data_out = 8'hFE;
                    16'h90EF: data_out = 8'hFF;
                    16'h90F0: data_out = 8'h80;
                    16'h90F1: data_out = 8'h81;
                    16'h90F2: data_out = 8'h82;
                    16'h90F3: data_out = 8'h83;
                    16'h90F4: data_out = 8'h84;
                    16'h90F5: data_out = 8'h85;
                    16'h90F6: data_out = 8'h86;
                    16'h90F7: data_out = 8'h87;
                    16'h90F8: data_out = 8'h88;
                    16'h90F9: data_out = 8'h89;
                    16'h90FA: data_out = 8'h8A;
                    16'h90FB: data_out = 8'h8B;
                    16'h90FC: data_out = 8'h8C;
                    16'h90FD: data_out = 8'h8D;
                    16'h90FE: data_out = 8'h8E;
                    16'h90FF: data_out = 8'h8F;
                    16'h9100: data_out = 8'h91;
                    16'h9101: data_out = 8'h90;
                    16'h9102: data_out = 8'h8F;
                    16'h9103: data_out = 8'h8E;
                    16'h9104: data_out = 8'h8D;
                    16'h9105: data_out = 8'h8C;
                    16'h9106: data_out = 8'h8B;
                    16'h9107: data_out = 8'h8A;
                    16'h9108: data_out = 8'h89;
                    16'h9109: data_out = 8'h88;
                    16'h910A: data_out = 8'h87;
                    16'h910B: data_out = 8'h86;
                    16'h910C: data_out = 8'h85;
                    16'h910D: data_out = 8'h84;
                    16'h910E: data_out = 8'h83;
                    16'h910F: data_out = 8'h82;
                    16'h9110: data_out = 8'h81;
                    16'h9111: data_out = 8'h0;
                    16'h9112: data_out = 8'h1;
                    16'h9113: data_out = 8'h2;
                    16'h9114: data_out = 8'h3;
                    16'h9115: data_out = 8'h4;
                    16'h9116: data_out = 8'h5;
                    16'h9117: data_out = 8'h6;
                    16'h9118: data_out = 8'h7;
                    16'h9119: data_out = 8'h8;
                    16'h911A: data_out = 8'h9;
                    16'h911B: data_out = 8'hA;
                    16'h911C: data_out = 8'hB;
                    16'h911D: data_out = 8'hC;
                    16'h911E: data_out = 8'hD;
                    16'h911F: data_out = 8'hE;
                    16'h9120: data_out = 8'hF;
                    16'h9121: data_out = 8'h10;
                    16'h9122: data_out = 8'h11;
                    16'h9123: data_out = 8'h12;
                    16'h9124: data_out = 8'h13;
                    16'h9125: data_out = 8'h14;
                    16'h9126: data_out = 8'h15;
                    16'h9127: data_out = 8'h16;
                    16'h9128: data_out = 8'h17;
                    16'h9129: data_out = 8'h18;
                    16'h912A: data_out = 8'h19;
                    16'h912B: data_out = 8'h1A;
                    16'h912C: data_out = 8'h1B;
                    16'h912D: data_out = 8'h1C;
                    16'h912E: data_out = 8'h1D;
                    16'h912F: data_out = 8'h1E;
                    16'h9130: data_out = 8'h1F;
                    16'h9131: data_out = 8'h20;
                    16'h9132: data_out = 8'h21;
                    16'h9133: data_out = 8'h22;
                    16'h9134: data_out = 8'h23;
                    16'h9135: data_out = 8'h24;
                    16'h9136: data_out = 8'h25;
                    16'h9137: data_out = 8'h26;
                    16'h9138: data_out = 8'h27;
                    16'h9139: data_out = 8'h28;
                    16'h913A: data_out = 8'h29;
                    16'h913B: data_out = 8'h2A;
                    16'h913C: data_out = 8'h2B;
                    16'h913D: data_out = 8'h2C;
                    16'h913E: data_out = 8'h2D;
                    16'h913F: data_out = 8'h2E;
                    16'h9140: data_out = 8'h2F;
                    16'h9141: data_out = 8'h30;
                    16'h9142: data_out = 8'h31;
                    16'h9143: data_out = 8'h32;
                    16'h9144: data_out = 8'h33;
                    16'h9145: data_out = 8'h34;
                    16'h9146: data_out = 8'h35;
                    16'h9147: data_out = 8'h36;
                    16'h9148: data_out = 8'h37;
                    16'h9149: data_out = 8'h38;
                    16'h914A: data_out = 8'h39;
                    16'h914B: data_out = 8'h3A;
                    16'h914C: data_out = 8'h3B;
                    16'h914D: data_out = 8'h3C;
                    16'h914E: data_out = 8'h3D;
                    16'h914F: data_out = 8'h3E;
                    16'h9150: data_out = 8'h3F;
                    16'h9151: data_out = 8'h40;
                    16'h9152: data_out = 8'h41;
                    16'h9153: data_out = 8'h42;
                    16'h9154: data_out = 8'h43;
                    16'h9155: data_out = 8'h44;
                    16'h9156: data_out = 8'h45;
                    16'h9157: data_out = 8'h46;
                    16'h9158: data_out = 8'h47;
                    16'h9159: data_out = 8'h48;
                    16'h915A: data_out = 8'h49;
                    16'h915B: data_out = 8'h4A;
                    16'h915C: data_out = 8'h4B;
                    16'h915D: data_out = 8'h4C;
                    16'h915E: data_out = 8'h4D;
                    16'h915F: data_out = 8'h4E;
                    16'h9160: data_out = 8'h4F;
                    16'h9161: data_out = 8'h50;
                    16'h9162: data_out = 8'h51;
                    16'h9163: data_out = 8'h52;
                    16'h9164: data_out = 8'h53;
                    16'h9165: data_out = 8'h54;
                    16'h9166: data_out = 8'h55;
                    16'h9167: data_out = 8'h56;
                    16'h9168: data_out = 8'h57;
                    16'h9169: data_out = 8'h58;
                    16'h916A: data_out = 8'h59;
                    16'h916B: data_out = 8'h5A;
                    16'h916C: data_out = 8'h5B;
                    16'h916D: data_out = 8'h5C;
                    16'h916E: data_out = 8'h5D;
                    16'h916F: data_out = 8'h5E;
                    16'h9170: data_out = 8'h5F;
                    16'h9171: data_out = 8'h60;
                    16'h9172: data_out = 8'h61;
                    16'h9173: data_out = 8'h62;
                    16'h9174: data_out = 8'h63;
                    16'h9175: data_out = 8'h64;
                    16'h9176: data_out = 8'h65;
                    16'h9177: data_out = 8'h66;
                    16'h9178: data_out = 8'h67;
                    16'h9179: data_out = 8'h68;
                    16'h917A: data_out = 8'h69;
                    16'h917B: data_out = 8'h6A;
                    16'h917C: data_out = 8'h6B;
                    16'h917D: data_out = 8'h6C;
                    16'h917E: data_out = 8'h6D;
                    16'h917F: data_out = 8'h6E;
                    16'h9180: data_out = 8'h91;
                    16'h9181: data_out = 8'h92;
                    16'h9182: data_out = 8'h93;
                    16'h9183: data_out = 8'h94;
                    16'h9184: data_out = 8'h95;
                    16'h9185: data_out = 8'h96;
                    16'h9186: data_out = 8'h97;
                    16'h9187: data_out = 8'h98;
                    16'h9188: data_out = 8'h99;
                    16'h9189: data_out = 8'h9A;
                    16'h918A: data_out = 8'h9B;
                    16'h918B: data_out = 8'h9C;
                    16'h918C: data_out = 8'h9D;
                    16'h918D: data_out = 8'h9E;
                    16'h918E: data_out = 8'h9F;
                    16'h918F: data_out = 8'hA0;
                    16'h9190: data_out = 8'hA1;
                    16'h9191: data_out = 8'hA2;
                    16'h9192: data_out = 8'hA3;
                    16'h9193: data_out = 8'hA4;
                    16'h9194: data_out = 8'hA5;
                    16'h9195: data_out = 8'hA6;
                    16'h9196: data_out = 8'hA7;
                    16'h9197: data_out = 8'hA8;
                    16'h9198: data_out = 8'hA9;
                    16'h9199: data_out = 8'hAA;
                    16'h919A: data_out = 8'hAB;
                    16'h919B: data_out = 8'hAC;
                    16'h919C: data_out = 8'hAD;
                    16'h919D: data_out = 8'hAE;
                    16'h919E: data_out = 8'hAF;
                    16'h919F: data_out = 8'hB0;
                    16'h91A0: data_out = 8'hB1;
                    16'h91A1: data_out = 8'hB2;
                    16'h91A2: data_out = 8'hB3;
                    16'h91A3: data_out = 8'hB4;
                    16'h91A4: data_out = 8'hB5;
                    16'h91A5: data_out = 8'hB6;
                    16'h91A6: data_out = 8'hB7;
                    16'h91A7: data_out = 8'hB8;
                    16'h91A8: data_out = 8'hB9;
                    16'h91A9: data_out = 8'hBA;
                    16'h91AA: data_out = 8'hBB;
                    16'h91AB: data_out = 8'hBC;
                    16'h91AC: data_out = 8'hBD;
                    16'h91AD: data_out = 8'hBE;
                    16'h91AE: data_out = 8'hBF;
                    16'h91AF: data_out = 8'hC0;
                    16'h91B0: data_out = 8'hC1;
                    16'h91B1: data_out = 8'hC2;
                    16'h91B2: data_out = 8'hC3;
                    16'h91B3: data_out = 8'hC4;
                    16'h91B4: data_out = 8'hC5;
                    16'h91B5: data_out = 8'hC6;
                    16'h91B6: data_out = 8'hC7;
                    16'h91B7: data_out = 8'hC8;
                    16'h91B8: data_out = 8'hC9;
                    16'h91B9: data_out = 8'hCA;
                    16'h91BA: data_out = 8'hCB;
                    16'h91BB: data_out = 8'hCC;
                    16'h91BC: data_out = 8'hCD;
                    16'h91BD: data_out = 8'hCE;
                    16'h91BE: data_out = 8'hCF;
                    16'h91BF: data_out = 8'hD0;
                    16'h91C0: data_out = 8'hD1;
                    16'h91C1: data_out = 8'hD2;
                    16'h91C2: data_out = 8'hD3;
                    16'h91C3: data_out = 8'hD4;
                    16'h91C4: data_out = 8'hD5;
                    16'h91C5: data_out = 8'hD6;
                    16'h91C6: data_out = 8'hD7;
                    16'h91C7: data_out = 8'hD8;
                    16'h91C8: data_out = 8'hD9;
                    16'h91C9: data_out = 8'hDA;
                    16'h91CA: data_out = 8'hDB;
                    16'h91CB: data_out = 8'hDC;
                    16'h91CC: data_out = 8'hDD;
                    16'h91CD: data_out = 8'hDE;
                    16'h91CE: data_out = 8'hDF;
                    16'h91CF: data_out = 8'hE0;
                    16'h91D0: data_out = 8'hE1;
                    16'h91D1: data_out = 8'hE2;
                    16'h91D2: data_out = 8'hE3;
                    16'h91D3: data_out = 8'hE4;
                    16'h91D4: data_out = 8'hE5;
                    16'h91D5: data_out = 8'hE6;
                    16'h91D6: data_out = 8'hE7;
                    16'h91D7: data_out = 8'hE8;
                    16'h91D8: data_out = 8'hE9;
                    16'h91D9: data_out = 8'hEA;
                    16'h91DA: data_out = 8'hEB;
                    16'h91DB: data_out = 8'hEC;
                    16'h91DC: data_out = 8'hED;
                    16'h91DD: data_out = 8'hEE;
                    16'h91DE: data_out = 8'hEF;
                    16'h91DF: data_out = 8'hF0;
                    16'h91E0: data_out = 8'hF1;
                    16'h91E1: data_out = 8'hF2;
                    16'h91E2: data_out = 8'hF3;
                    16'h91E3: data_out = 8'hF4;
                    16'h91E4: data_out = 8'hF5;
                    16'h91E5: data_out = 8'hF6;
                    16'h91E6: data_out = 8'hF7;
                    16'h91E7: data_out = 8'hF8;
                    16'h91E8: data_out = 8'hF9;
                    16'h91E9: data_out = 8'hFA;
                    16'h91EA: data_out = 8'hFB;
                    16'h91EB: data_out = 8'hFC;
                    16'h91EC: data_out = 8'hFD;
                    16'h91ED: data_out = 8'hFE;
                    16'h91EE: data_out = 8'hFF;
                    16'h91EF: data_out = 8'h80;
                    16'h91F0: data_out = 8'h81;
                    16'h91F1: data_out = 8'h82;
                    16'h91F2: data_out = 8'h83;
                    16'h91F3: data_out = 8'h84;
                    16'h91F4: data_out = 8'h85;
                    16'h91F5: data_out = 8'h86;
                    16'h91F6: data_out = 8'h87;
                    16'h91F7: data_out = 8'h88;
                    16'h91F8: data_out = 8'h89;
                    16'h91F9: data_out = 8'h8A;
                    16'h91FA: data_out = 8'h8B;
                    16'h91FB: data_out = 8'h8C;
                    16'h91FC: data_out = 8'h8D;
                    16'h91FD: data_out = 8'h8E;
                    16'h91FE: data_out = 8'h8F;
                    16'h91FF: data_out = 8'h90;
                    16'h9200: data_out = 8'h92;
                    16'h9201: data_out = 8'h91;
                    16'h9202: data_out = 8'h90;
                    16'h9203: data_out = 8'h8F;
                    16'h9204: data_out = 8'h8E;
                    16'h9205: data_out = 8'h8D;
                    16'h9206: data_out = 8'h8C;
                    16'h9207: data_out = 8'h8B;
                    16'h9208: data_out = 8'h8A;
                    16'h9209: data_out = 8'h89;
                    16'h920A: data_out = 8'h88;
                    16'h920B: data_out = 8'h87;
                    16'h920C: data_out = 8'h86;
                    16'h920D: data_out = 8'h85;
                    16'h920E: data_out = 8'h84;
                    16'h920F: data_out = 8'h83;
                    16'h9210: data_out = 8'h82;
                    16'h9211: data_out = 8'h81;
                    16'h9212: data_out = 8'h0;
                    16'h9213: data_out = 8'h1;
                    16'h9214: data_out = 8'h2;
                    16'h9215: data_out = 8'h3;
                    16'h9216: data_out = 8'h4;
                    16'h9217: data_out = 8'h5;
                    16'h9218: data_out = 8'h6;
                    16'h9219: data_out = 8'h7;
                    16'h921A: data_out = 8'h8;
                    16'h921B: data_out = 8'h9;
                    16'h921C: data_out = 8'hA;
                    16'h921D: data_out = 8'hB;
                    16'h921E: data_out = 8'hC;
                    16'h921F: data_out = 8'hD;
                    16'h9220: data_out = 8'hE;
                    16'h9221: data_out = 8'hF;
                    16'h9222: data_out = 8'h10;
                    16'h9223: data_out = 8'h11;
                    16'h9224: data_out = 8'h12;
                    16'h9225: data_out = 8'h13;
                    16'h9226: data_out = 8'h14;
                    16'h9227: data_out = 8'h15;
                    16'h9228: data_out = 8'h16;
                    16'h9229: data_out = 8'h17;
                    16'h922A: data_out = 8'h18;
                    16'h922B: data_out = 8'h19;
                    16'h922C: data_out = 8'h1A;
                    16'h922D: data_out = 8'h1B;
                    16'h922E: data_out = 8'h1C;
                    16'h922F: data_out = 8'h1D;
                    16'h9230: data_out = 8'h1E;
                    16'h9231: data_out = 8'h1F;
                    16'h9232: data_out = 8'h20;
                    16'h9233: data_out = 8'h21;
                    16'h9234: data_out = 8'h22;
                    16'h9235: data_out = 8'h23;
                    16'h9236: data_out = 8'h24;
                    16'h9237: data_out = 8'h25;
                    16'h9238: data_out = 8'h26;
                    16'h9239: data_out = 8'h27;
                    16'h923A: data_out = 8'h28;
                    16'h923B: data_out = 8'h29;
                    16'h923C: data_out = 8'h2A;
                    16'h923D: data_out = 8'h2B;
                    16'h923E: data_out = 8'h2C;
                    16'h923F: data_out = 8'h2D;
                    16'h9240: data_out = 8'h2E;
                    16'h9241: data_out = 8'h2F;
                    16'h9242: data_out = 8'h30;
                    16'h9243: data_out = 8'h31;
                    16'h9244: data_out = 8'h32;
                    16'h9245: data_out = 8'h33;
                    16'h9246: data_out = 8'h34;
                    16'h9247: data_out = 8'h35;
                    16'h9248: data_out = 8'h36;
                    16'h9249: data_out = 8'h37;
                    16'h924A: data_out = 8'h38;
                    16'h924B: data_out = 8'h39;
                    16'h924C: data_out = 8'h3A;
                    16'h924D: data_out = 8'h3B;
                    16'h924E: data_out = 8'h3C;
                    16'h924F: data_out = 8'h3D;
                    16'h9250: data_out = 8'h3E;
                    16'h9251: data_out = 8'h3F;
                    16'h9252: data_out = 8'h40;
                    16'h9253: data_out = 8'h41;
                    16'h9254: data_out = 8'h42;
                    16'h9255: data_out = 8'h43;
                    16'h9256: data_out = 8'h44;
                    16'h9257: data_out = 8'h45;
                    16'h9258: data_out = 8'h46;
                    16'h9259: data_out = 8'h47;
                    16'h925A: data_out = 8'h48;
                    16'h925B: data_out = 8'h49;
                    16'h925C: data_out = 8'h4A;
                    16'h925D: data_out = 8'h4B;
                    16'h925E: data_out = 8'h4C;
                    16'h925F: data_out = 8'h4D;
                    16'h9260: data_out = 8'h4E;
                    16'h9261: data_out = 8'h4F;
                    16'h9262: data_out = 8'h50;
                    16'h9263: data_out = 8'h51;
                    16'h9264: data_out = 8'h52;
                    16'h9265: data_out = 8'h53;
                    16'h9266: data_out = 8'h54;
                    16'h9267: data_out = 8'h55;
                    16'h9268: data_out = 8'h56;
                    16'h9269: data_out = 8'h57;
                    16'h926A: data_out = 8'h58;
                    16'h926B: data_out = 8'h59;
                    16'h926C: data_out = 8'h5A;
                    16'h926D: data_out = 8'h5B;
                    16'h926E: data_out = 8'h5C;
                    16'h926F: data_out = 8'h5D;
                    16'h9270: data_out = 8'h5E;
                    16'h9271: data_out = 8'h5F;
                    16'h9272: data_out = 8'h60;
                    16'h9273: data_out = 8'h61;
                    16'h9274: data_out = 8'h62;
                    16'h9275: data_out = 8'h63;
                    16'h9276: data_out = 8'h64;
                    16'h9277: data_out = 8'h65;
                    16'h9278: data_out = 8'h66;
                    16'h9279: data_out = 8'h67;
                    16'h927A: data_out = 8'h68;
                    16'h927B: data_out = 8'h69;
                    16'h927C: data_out = 8'h6A;
                    16'h927D: data_out = 8'h6B;
                    16'h927E: data_out = 8'h6C;
                    16'h927F: data_out = 8'h6D;
                    16'h9280: data_out = 8'h92;
                    16'h9281: data_out = 8'h93;
                    16'h9282: data_out = 8'h94;
                    16'h9283: data_out = 8'h95;
                    16'h9284: data_out = 8'h96;
                    16'h9285: data_out = 8'h97;
                    16'h9286: data_out = 8'h98;
                    16'h9287: data_out = 8'h99;
                    16'h9288: data_out = 8'h9A;
                    16'h9289: data_out = 8'h9B;
                    16'h928A: data_out = 8'h9C;
                    16'h928B: data_out = 8'h9D;
                    16'h928C: data_out = 8'h9E;
                    16'h928D: data_out = 8'h9F;
                    16'h928E: data_out = 8'hA0;
                    16'h928F: data_out = 8'hA1;
                    16'h9290: data_out = 8'hA2;
                    16'h9291: data_out = 8'hA3;
                    16'h9292: data_out = 8'hA4;
                    16'h9293: data_out = 8'hA5;
                    16'h9294: data_out = 8'hA6;
                    16'h9295: data_out = 8'hA7;
                    16'h9296: data_out = 8'hA8;
                    16'h9297: data_out = 8'hA9;
                    16'h9298: data_out = 8'hAA;
                    16'h9299: data_out = 8'hAB;
                    16'h929A: data_out = 8'hAC;
                    16'h929B: data_out = 8'hAD;
                    16'h929C: data_out = 8'hAE;
                    16'h929D: data_out = 8'hAF;
                    16'h929E: data_out = 8'hB0;
                    16'h929F: data_out = 8'hB1;
                    16'h92A0: data_out = 8'hB2;
                    16'h92A1: data_out = 8'hB3;
                    16'h92A2: data_out = 8'hB4;
                    16'h92A3: data_out = 8'hB5;
                    16'h92A4: data_out = 8'hB6;
                    16'h92A5: data_out = 8'hB7;
                    16'h92A6: data_out = 8'hB8;
                    16'h92A7: data_out = 8'hB9;
                    16'h92A8: data_out = 8'hBA;
                    16'h92A9: data_out = 8'hBB;
                    16'h92AA: data_out = 8'hBC;
                    16'h92AB: data_out = 8'hBD;
                    16'h92AC: data_out = 8'hBE;
                    16'h92AD: data_out = 8'hBF;
                    16'h92AE: data_out = 8'hC0;
                    16'h92AF: data_out = 8'hC1;
                    16'h92B0: data_out = 8'hC2;
                    16'h92B1: data_out = 8'hC3;
                    16'h92B2: data_out = 8'hC4;
                    16'h92B3: data_out = 8'hC5;
                    16'h92B4: data_out = 8'hC6;
                    16'h92B5: data_out = 8'hC7;
                    16'h92B6: data_out = 8'hC8;
                    16'h92B7: data_out = 8'hC9;
                    16'h92B8: data_out = 8'hCA;
                    16'h92B9: data_out = 8'hCB;
                    16'h92BA: data_out = 8'hCC;
                    16'h92BB: data_out = 8'hCD;
                    16'h92BC: data_out = 8'hCE;
                    16'h92BD: data_out = 8'hCF;
                    16'h92BE: data_out = 8'hD0;
                    16'h92BF: data_out = 8'hD1;
                    16'h92C0: data_out = 8'hD2;
                    16'h92C1: data_out = 8'hD3;
                    16'h92C2: data_out = 8'hD4;
                    16'h92C3: data_out = 8'hD5;
                    16'h92C4: data_out = 8'hD6;
                    16'h92C5: data_out = 8'hD7;
                    16'h92C6: data_out = 8'hD8;
                    16'h92C7: data_out = 8'hD9;
                    16'h92C8: data_out = 8'hDA;
                    16'h92C9: data_out = 8'hDB;
                    16'h92CA: data_out = 8'hDC;
                    16'h92CB: data_out = 8'hDD;
                    16'h92CC: data_out = 8'hDE;
                    16'h92CD: data_out = 8'hDF;
                    16'h92CE: data_out = 8'hE0;
                    16'h92CF: data_out = 8'hE1;
                    16'h92D0: data_out = 8'hE2;
                    16'h92D1: data_out = 8'hE3;
                    16'h92D2: data_out = 8'hE4;
                    16'h92D3: data_out = 8'hE5;
                    16'h92D4: data_out = 8'hE6;
                    16'h92D5: data_out = 8'hE7;
                    16'h92D6: data_out = 8'hE8;
                    16'h92D7: data_out = 8'hE9;
                    16'h92D8: data_out = 8'hEA;
                    16'h92D9: data_out = 8'hEB;
                    16'h92DA: data_out = 8'hEC;
                    16'h92DB: data_out = 8'hED;
                    16'h92DC: data_out = 8'hEE;
                    16'h92DD: data_out = 8'hEF;
                    16'h92DE: data_out = 8'hF0;
                    16'h92DF: data_out = 8'hF1;
                    16'h92E0: data_out = 8'hF2;
                    16'h92E1: data_out = 8'hF3;
                    16'h92E2: data_out = 8'hF4;
                    16'h92E3: data_out = 8'hF5;
                    16'h92E4: data_out = 8'hF6;
                    16'h92E5: data_out = 8'hF7;
                    16'h92E6: data_out = 8'hF8;
                    16'h92E7: data_out = 8'hF9;
                    16'h92E8: data_out = 8'hFA;
                    16'h92E9: data_out = 8'hFB;
                    16'h92EA: data_out = 8'hFC;
                    16'h92EB: data_out = 8'hFD;
                    16'h92EC: data_out = 8'hFE;
                    16'h92ED: data_out = 8'hFF;
                    16'h92EE: data_out = 8'h80;
                    16'h92EF: data_out = 8'h81;
                    16'h92F0: data_out = 8'h82;
                    16'h92F1: data_out = 8'h83;
                    16'h92F2: data_out = 8'h84;
                    16'h92F3: data_out = 8'h85;
                    16'h92F4: data_out = 8'h86;
                    16'h92F5: data_out = 8'h87;
                    16'h92F6: data_out = 8'h88;
                    16'h92F7: data_out = 8'h89;
                    16'h92F8: data_out = 8'h8A;
                    16'h92F9: data_out = 8'h8B;
                    16'h92FA: data_out = 8'h8C;
                    16'h92FB: data_out = 8'h8D;
                    16'h92FC: data_out = 8'h8E;
                    16'h92FD: data_out = 8'h8F;
                    16'h92FE: data_out = 8'h90;
                    16'h92FF: data_out = 8'h91;
                    16'h9300: data_out = 8'h93;
                    16'h9301: data_out = 8'h92;
                    16'h9302: data_out = 8'h91;
                    16'h9303: data_out = 8'h90;
                    16'h9304: data_out = 8'h8F;
                    16'h9305: data_out = 8'h8E;
                    16'h9306: data_out = 8'h8D;
                    16'h9307: data_out = 8'h8C;
                    16'h9308: data_out = 8'h8B;
                    16'h9309: data_out = 8'h8A;
                    16'h930A: data_out = 8'h89;
                    16'h930B: data_out = 8'h88;
                    16'h930C: data_out = 8'h87;
                    16'h930D: data_out = 8'h86;
                    16'h930E: data_out = 8'h85;
                    16'h930F: data_out = 8'h84;
                    16'h9310: data_out = 8'h83;
                    16'h9311: data_out = 8'h82;
                    16'h9312: data_out = 8'h81;
                    16'h9313: data_out = 8'h0;
                    16'h9314: data_out = 8'h1;
                    16'h9315: data_out = 8'h2;
                    16'h9316: data_out = 8'h3;
                    16'h9317: data_out = 8'h4;
                    16'h9318: data_out = 8'h5;
                    16'h9319: data_out = 8'h6;
                    16'h931A: data_out = 8'h7;
                    16'h931B: data_out = 8'h8;
                    16'h931C: data_out = 8'h9;
                    16'h931D: data_out = 8'hA;
                    16'h931E: data_out = 8'hB;
                    16'h931F: data_out = 8'hC;
                    16'h9320: data_out = 8'hD;
                    16'h9321: data_out = 8'hE;
                    16'h9322: data_out = 8'hF;
                    16'h9323: data_out = 8'h10;
                    16'h9324: data_out = 8'h11;
                    16'h9325: data_out = 8'h12;
                    16'h9326: data_out = 8'h13;
                    16'h9327: data_out = 8'h14;
                    16'h9328: data_out = 8'h15;
                    16'h9329: data_out = 8'h16;
                    16'h932A: data_out = 8'h17;
                    16'h932B: data_out = 8'h18;
                    16'h932C: data_out = 8'h19;
                    16'h932D: data_out = 8'h1A;
                    16'h932E: data_out = 8'h1B;
                    16'h932F: data_out = 8'h1C;
                    16'h9330: data_out = 8'h1D;
                    16'h9331: data_out = 8'h1E;
                    16'h9332: data_out = 8'h1F;
                    16'h9333: data_out = 8'h20;
                    16'h9334: data_out = 8'h21;
                    16'h9335: data_out = 8'h22;
                    16'h9336: data_out = 8'h23;
                    16'h9337: data_out = 8'h24;
                    16'h9338: data_out = 8'h25;
                    16'h9339: data_out = 8'h26;
                    16'h933A: data_out = 8'h27;
                    16'h933B: data_out = 8'h28;
                    16'h933C: data_out = 8'h29;
                    16'h933D: data_out = 8'h2A;
                    16'h933E: data_out = 8'h2B;
                    16'h933F: data_out = 8'h2C;
                    16'h9340: data_out = 8'h2D;
                    16'h9341: data_out = 8'h2E;
                    16'h9342: data_out = 8'h2F;
                    16'h9343: data_out = 8'h30;
                    16'h9344: data_out = 8'h31;
                    16'h9345: data_out = 8'h32;
                    16'h9346: data_out = 8'h33;
                    16'h9347: data_out = 8'h34;
                    16'h9348: data_out = 8'h35;
                    16'h9349: data_out = 8'h36;
                    16'h934A: data_out = 8'h37;
                    16'h934B: data_out = 8'h38;
                    16'h934C: data_out = 8'h39;
                    16'h934D: data_out = 8'h3A;
                    16'h934E: data_out = 8'h3B;
                    16'h934F: data_out = 8'h3C;
                    16'h9350: data_out = 8'h3D;
                    16'h9351: data_out = 8'h3E;
                    16'h9352: data_out = 8'h3F;
                    16'h9353: data_out = 8'h40;
                    16'h9354: data_out = 8'h41;
                    16'h9355: data_out = 8'h42;
                    16'h9356: data_out = 8'h43;
                    16'h9357: data_out = 8'h44;
                    16'h9358: data_out = 8'h45;
                    16'h9359: data_out = 8'h46;
                    16'h935A: data_out = 8'h47;
                    16'h935B: data_out = 8'h48;
                    16'h935C: data_out = 8'h49;
                    16'h935D: data_out = 8'h4A;
                    16'h935E: data_out = 8'h4B;
                    16'h935F: data_out = 8'h4C;
                    16'h9360: data_out = 8'h4D;
                    16'h9361: data_out = 8'h4E;
                    16'h9362: data_out = 8'h4F;
                    16'h9363: data_out = 8'h50;
                    16'h9364: data_out = 8'h51;
                    16'h9365: data_out = 8'h52;
                    16'h9366: data_out = 8'h53;
                    16'h9367: data_out = 8'h54;
                    16'h9368: data_out = 8'h55;
                    16'h9369: data_out = 8'h56;
                    16'h936A: data_out = 8'h57;
                    16'h936B: data_out = 8'h58;
                    16'h936C: data_out = 8'h59;
                    16'h936D: data_out = 8'h5A;
                    16'h936E: data_out = 8'h5B;
                    16'h936F: data_out = 8'h5C;
                    16'h9370: data_out = 8'h5D;
                    16'h9371: data_out = 8'h5E;
                    16'h9372: data_out = 8'h5F;
                    16'h9373: data_out = 8'h60;
                    16'h9374: data_out = 8'h61;
                    16'h9375: data_out = 8'h62;
                    16'h9376: data_out = 8'h63;
                    16'h9377: data_out = 8'h64;
                    16'h9378: data_out = 8'h65;
                    16'h9379: data_out = 8'h66;
                    16'h937A: data_out = 8'h67;
                    16'h937B: data_out = 8'h68;
                    16'h937C: data_out = 8'h69;
                    16'h937D: data_out = 8'h6A;
                    16'h937E: data_out = 8'h6B;
                    16'h937F: data_out = 8'h6C;
                    16'h9380: data_out = 8'h93;
                    16'h9381: data_out = 8'h94;
                    16'h9382: data_out = 8'h95;
                    16'h9383: data_out = 8'h96;
                    16'h9384: data_out = 8'h97;
                    16'h9385: data_out = 8'h98;
                    16'h9386: data_out = 8'h99;
                    16'h9387: data_out = 8'h9A;
                    16'h9388: data_out = 8'h9B;
                    16'h9389: data_out = 8'h9C;
                    16'h938A: data_out = 8'h9D;
                    16'h938B: data_out = 8'h9E;
                    16'h938C: data_out = 8'h9F;
                    16'h938D: data_out = 8'hA0;
                    16'h938E: data_out = 8'hA1;
                    16'h938F: data_out = 8'hA2;
                    16'h9390: data_out = 8'hA3;
                    16'h9391: data_out = 8'hA4;
                    16'h9392: data_out = 8'hA5;
                    16'h9393: data_out = 8'hA6;
                    16'h9394: data_out = 8'hA7;
                    16'h9395: data_out = 8'hA8;
                    16'h9396: data_out = 8'hA9;
                    16'h9397: data_out = 8'hAA;
                    16'h9398: data_out = 8'hAB;
                    16'h9399: data_out = 8'hAC;
                    16'h939A: data_out = 8'hAD;
                    16'h939B: data_out = 8'hAE;
                    16'h939C: data_out = 8'hAF;
                    16'h939D: data_out = 8'hB0;
                    16'h939E: data_out = 8'hB1;
                    16'h939F: data_out = 8'hB2;
                    16'h93A0: data_out = 8'hB3;
                    16'h93A1: data_out = 8'hB4;
                    16'h93A2: data_out = 8'hB5;
                    16'h93A3: data_out = 8'hB6;
                    16'h93A4: data_out = 8'hB7;
                    16'h93A5: data_out = 8'hB8;
                    16'h93A6: data_out = 8'hB9;
                    16'h93A7: data_out = 8'hBA;
                    16'h93A8: data_out = 8'hBB;
                    16'h93A9: data_out = 8'hBC;
                    16'h93AA: data_out = 8'hBD;
                    16'h93AB: data_out = 8'hBE;
                    16'h93AC: data_out = 8'hBF;
                    16'h93AD: data_out = 8'hC0;
                    16'h93AE: data_out = 8'hC1;
                    16'h93AF: data_out = 8'hC2;
                    16'h93B0: data_out = 8'hC3;
                    16'h93B1: data_out = 8'hC4;
                    16'h93B2: data_out = 8'hC5;
                    16'h93B3: data_out = 8'hC6;
                    16'h93B4: data_out = 8'hC7;
                    16'h93B5: data_out = 8'hC8;
                    16'h93B6: data_out = 8'hC9;
                    16'h93B7: data_out = 8'hCA;
                    16'h93B8: data_out = 8'hCB;
                    16'h93B9: data_out = 8'hCC;
                    16'h93BA: data_out = 8'hCD;
                    16'h93BB: data_out = 8'hCE;
                    16'h93BC: data_out = 8'hCF;
                    16'h93BD: data_out = 8'hD0;
                    16'h93BE: data_out = 8'hD1;
                    16'h93BF: data_out = 8'hD2;
                    16'h93C0: data_out = 8'hD3;
                    16'h93C1: data_out = 8'hD4;
                    16'h93C2: data_out = 8'hD5;
                    16'h93C3: data_out = 8'hD6;
                    16'h93C4: data_out = 8'hD7;
                    16'h93C5: data_out = 8'hD8;
                    16'h93C6: data_out = 8'hD9;
                    16'h93C7: data_out = 8'hDA;
                    16'h93C8: data_out = 8'hDB;
                    16'h93C9: data_out = 8'hDC;
                    16'h93CA: data_out = 8'hDD;
                    16'h93CB: data_out = 8'hDE;
                    16'h93CC: data_out = 8'hDF;
                    16'h93CD: data_out = 8'hE0;
                    16'h93CE: data_out = 8'hE1;
                    16'h93CF: data_out = 8'hE2;
                    16'h93D0: data_out = 8'hE3;
                    16'h93D1: data_out = 8'hE4;
                    16'h93D2: data_out = 8'hE5;
                    16'h93D3: data_out = 8'hE6;
                    16'h93D4: data_out = 8'hE7;
                    16'h93D5: data_out = 8'hE8;
                    16'h93D6: data_out = 8'hE9;
                    16'h93D7: data_out = 8'hEA;
                    16'h93D8: data_out = 8'hEB;
                    16'h93D9: data_out = 8'hEC;
                    16'h93DA: data_out = 8'hED;
                    16'h93DB: data_out = 8'hEE;
                    16'h93DC: data_out = 8'hEF;
                    16'h93DD: data_out = 8'hF0;
                    16'h93DE: data_out = 8'hF1;
                    16'h93DF: data_out = 8'hF2;
                    16'h93E0: data_out = 8'hF3;
                    16'h93E1: data_out = 8'hF4;
                    16'h93E2: data_out = 8'hF5;
                    16'h93E3: data_out = 8'hF6;
                    16'h93E4: data_out = 8'hF7;
                    16'h93E5: data_out = 8'hF8;
                    16'h93E6: data_out = 8'hF9;
                    16'h93E7: data_out = 8'hFA;
                    16'h93E8: data_out = 8'hFB;
                    16'h93E9: data_out = 8'hFC;
                    16'h93EA: data_out = 8'hFD;
                    16'h93EB: data_out = 8'hFE;
                    16'h93EC: data_out = 8'hFF;
                    16'h93ED: data_out = 8'h80;
                    16'h93EE: data_out = 8'h81;
                    16'h93EF: data_out = 8'h82;
                    16'h93F0: data_out = 8'h83;
                    16'h93F1: data_out = 8'h84;
                    16'h93F2: data_out = 8'h85;
                    16'h93F3: data_out = 8'h86;
                    16'h93F4: data_out = 8'h87;
                    16'h93F5: data_out = 8'h88;
                    16'h93F6: data_out = 8'h89;
                    16'h93F7: data_out = 8'h8A;
                    16'h93F8: data_out = 8'h8B;
                    16'h93F9: data_out = 8'h8C;
                    16'h93FA: data_out = 8'h8D;
                    16'h93FB: data_out = 8'h8E;
                    16'h93FC: data_out = 8'h8F;
                    16'h93FD: data_out = 8'h90;
                    16'h93FE: data_out = 8'h91;
                    16'h93FF: data_out = 8'h92;
                    16'h9400: data_out = 8'h94;
                    16'h9401: data_out = 8'h93;
                    16'h9402: data_out = 8'h92;
                    16'h9403: data_out = 8'h91;
                    16'h9404: data_out = 8'h90;
                    16'h9405: data_out = 8'h8F;
                    16'h9406: data_out = 8'h8E;
                    16'h9407: data_out = 8'h8D;
                    16'h9408: data_out = 8'h8C;
                    16'h9409: data_out = 8'h8B;
                    16'h940A: data_out = 8'h8A;
                    16'h940B: data_out = 8'h89;
                    16'h940C: data_out = 8'h88;
                    16'h940D: data_out = 8'h87;
                    16'h940E: data_out = 8'h86;
                    16'h940F: data_out = 8'h85;
                    16'h9410: data_out = 8'h84;
                    16'h9411: data_out = 8'h83;
                    16'h9412: data_out = 8'h82;
                    16'h9413: data_out = 8'h81;
                    16'h9414: data_out = 8'h0;
                    16'h9415: data_out = 8'h1;
                    16'h9416: data_out = 8'h2;
                    16'h9417: data_out = 8'h3;
                    16'h9418: data_out = 8'h4;
                    16'h9419: data_out = 8'h5;
                    16'h941A: data_out = 8'h6;
                    16'h941B: data_out = 8'h7;
                    16'h941C: data_out = 8'h8;
                    16'h941D: data_out = 8'h9;
                    16'h941E: data_out = 8'hA;
                    16'h941F: data_out = 8'hB;
                    16'h9420: data_out = 8'hC;
                    16'h9421: data_out = 8'hD;
                    16'h9422: data_out = 8'hE;
                    16'h9423: data_out = 8'hF;
                    16'h9424: data_out = 8'h10;
                    16'h9425: data_out = 8'h11;
                    16'h9426: data_out = 8'h12;
                    16'h9427: data_out = 8'h13;
                    16'h9428: data_out = 8'h14;
                    16'h9429: data_out = 8'h15;
                    16'h942A: data_out = 8'h16;
                    16'h942B: data_out = 8'h17;
                    16'h942C: data_out = 8'h18;
                    16'h942D: data_out = 8'h19;
                    16'h942E: data_out = 8'h1A;
                    16'h942F: data_out = 8'h1B;
                    16'h9430: data_out = 8'h1C;
                    16'h9431: data_out = 8'h1D;
                    16'h9432: data_out = 8'h1E;
                    16'h9433: data_out = 8'h1F;
                    16'h9434: data_out = 8'h20;
                    16'h9435: data_out = 8'h21;
                    16'h9436: data_out = 8'h22;
                    16'h9437: data_out = 8'h23;
                    16'h9438: data_out = 8'h24;
                    16'h9439: data_out = 8'h25;
                    16'h943A: data_out = 8'h26;
                    16'h943B: data_out = 8'h27;
                    16'h943C: data_out = 8'h28;
                    16'h943D: data_out = 8'h29;
                    16'h943E: data_out = 8'h2A;
                    16'h943F: data_out = 8'h2B;
                    16'h9440: data_out = 8'h2C;
                    16'h9441: data_out = 8'h2D;
                    16'h9442: data_out = 8'h2E;
                    16'h9443: data_out = 8'h2F;
                    16'h9444: data_out = 8'h30;
                    16'h9445: data_out = 8'h31;
                    16'h9446: data_out = 8'h32;
                    16'h9447: data_out = 8'h33;
                    16'h9448: data_out = 8'h34;
                    16'h9449: data_out = 8'h35;
                    16'h944A: data_out = 8'h36;
                    16'h944B: data_out = 8'h37;
                    16'h944C: data_out = 8'h38;
                    16'h944D: data_out = 8'h39;
                    16'h944E: data_out = 8'h3A;
                    16'h944F: data_out = 8'h3B;
                    16'h9450: data_out = 8'h3C;
                    16'h9451: data_out = 8'h3D;
                    16'h9452: data_out = 8'h3E;
                    16'h9453: data_out = 8'h3F;
                    16'h9454: data_out = 8'h40;
                    16'h9455: data_out = 8'h41;
                    16'h9456: data_out = 8'h42;
                    16'h9457: data_out = 8'h43;
                    16'h9458: data_out = 8'h44;
                    16'h9459: data_out = 8'h45;
                    16'h945A: data_out = 8'h46;
                    16'h945B: data_out = 8'h47;
                    16'h945C: data_out = 8'h48;
                    16'h945D: data_out = 8'h49;
                    16'h945E: data_out = 8'h4A;
                    16'h945F: data_out = 8'h4B;
                    16'h9460: data_out = 8'h4C;
                    16'h9461: data_out = 8'h4D;
                    16'h9462: data_out = 8'h4E;
                    16'h9463: data_out = 8'h4F;
                    16'h9464: data_out = 8'h50;
                    16'h9465: data_out = 8'h51;
                    16'h9466: data_out = 8'h52;
                    16'h9467: data_out = 8'h53;
                    16'h9468: data_out = 8'h54;
                    16'h9469: data_out = 8'h55;
                    16'h946A: data_out = 8'h56;
                    16'h946B: data_out = 8'h57;
                    16'h946C: data_out = 8'h58;
                    16'h946D: data_out = 8'h59;
                    16'h946E: data_out = 8'h5A;
                    16'h946F: data_out = 8'h5B;
                    16'h9470: data_out = 8'h5C;
                    16'h9471: data_out = 8'h5D;
                    16'h9472: data_out = 8'h5E;
                    16'h9473: data_out = 8'h5F;
                    16'h9474: data_out = 8'h60;
                    16'h9475: data_out = 8'h61;
                    16'h9476: data_out = 8'h62;
                    16'h9477: data_out = 8'h63;
                    16'h9478: data_out = 8'h64;
                    16'h9479: data_out = 8'h65;
                    16'h947A: data_out = 8'h66;
                    16'h947B: data_out = 8'h67;
                    16'h947C: data_out = 8'h68;
                    16'h947D: data_out = 8'h69;
                    16'h947E: data_out = 8'h6A;
                    16'h947F: data_out = 8'h6B;
                    16'h9480: data_out = 8'h94;
                    16'h9481: data_out = 8'h95;
                    16'h9482: data_out = 8'h96;
                    16'h9483: data_out = 8'h97;
                    16'h9484: data_out = 8'h98;
                    16'h9485: data_out = 8'h99;
                    16'h9486: data_out = 8'h9A;
                    16'h9487: data_out = 8'h9B;
                    16'h9488: data_out = 8'h9C;
                    16'h9489: data_out = 8'h9D;
                    16'h948A: data_out = 8'h9E;
                    16'h948B: data_out = 8'h9F;
                    16'h948C: data_out = 8'hA0;
                    16'h948D: data_out = 8'hA1;
                    16'h948E: data_out = 8'hA2;
                    16'h948F: data_out = 8'hA3;
                    16'h9490: data_out = 8'hA4;
                    16'h9491: data_out = 8'hA5;
                    16'h9492: data_out = 8'hA6;
                    16'h9493: data_out = 8'hA7;
                    16'h9494: data_out = 8'hA8;
                    16'h9495: data_out = 8'hA9;
                    16'h9496: data_out = 8'hAA;
                    16'h9497: data_out = 8'hAB;
                    16'h9498: data_out = 8'hAC;
                    16'h9499: data_out = 8'hAD;
                    16'h949A: data_out = 8'hAE;
                    16'h949B: data_out = 8'hAF;
                    16'h949C: data_out = 8'hB0;
                    16'h949D: data_out = 8'hB1;
                    16'h949E: data_out = 8'hB2;
                    16'h949F: data_out = 8'hB3;
                    16'h94A0: data_out = 8'hB4;
                    16'h94A1: data_out = 8'hB5;
                    16'h94A2: data_out = 8'hB6;
                    16'h94A3: data_out = 8'hB7;
                    16'h94A4: data_out = 8'hB8;
                    16'h94A5: data_out = 8'hB9;
                    16'h94A6: data_out = 8'hBA;
                    16'h94A7: data_out = 8'hBB;
                    16'h94A8: data_out = 8'hBC;
                    16'h94A9: data_out = 8'hBD;
                    16'h94AA: data_out = 8'hBE;
                    16'h94AB: data_out = 8'hBF;
                    16'h94AC: data_out = 8'hC0;
                    16'h94AD: data_out = 8'hC1;
                    16'h94AE: data_out = 8'hC2;
                    16'h94AF: data_out = 8'hC3;
                    16'h94B0: data_out = 8'hC4;
                    16'h94B1: data_out = 8'hC5;
                    16'h94B2: data_out = 8'hC6;
                    16'h94B3: data_out = 8'hC7;
                    16'h94B4: data_out = 8'hC8;
                    16'h94B5: data_out = 8'hC9;
                    16'h94B6: data_out = 8'hCA;
                    16'h94B7: data_out = 8'hCB;
                    16'h94B8: data_out = 8'hCC;
                    16'h94B9: data_out = 8'hCD;
                    16'h94BA: data_out = 8'hCE;
                    16'h94BB: data_out = 8'hCF;
                    16'h94BC: data_out = 8'hD0;
                    16'h94BD: data_out = 8'hD1;
                    16'h94BE: data_out = 8'hD2;
                    16'h94BF: data_out = 8'hD3;
                    16'h94C0: data_out = 8'hD4;
                    16'h94C1: data_out = 8'hD5;
                    16'h94C2: data_out = 8'hD6;
                    16'h94C3: data_out = 8'hD7;
                    16'h94C4: data_out = 8'hD8;
                    16'h94C5: data_out = 8'hD9;
                    16'h94C6: data_out = 8'hDA;
                    16'h94C7: data_out = 8'hDB;
                    16'h94C8: data_out = 8'hDC;
                    16'h94C9: data_out = 8'hDD;
                    16'h94CA: data_out = 8'hDE;
                    16'h94CB: data_out = 8'hDF;
                    16'h94CC: data_out = 8'hE0;
                    16'h94CD: data_out = 8'hE1;
                    16'h94CE: data_out = 8'hE2;
                    16'h94CF: data_out = 8'hE3;
                    16'h94D0: data_out = 8'hE4;
                    16'h94D1: data_out = 8'hE5;
                    16'h94D2: data_out = 8'hE6;
                    16'h94D3: data_out = 8'hE7;
                    16'h94D4: data_out = 8'hE8;
                    16'h94D5: data_out = 8'hE9;
                    16'h94D6: data_out = 8'hEA;
                    16'h94D7: data_out = 8'hEB;
                    16'h94D8: data_out = 8'hEC;
                    16'h94D9: data_out = 8'hED;
                    16'h94DA: data_out = 8'hEE;
                    16'h94DB: data_out = 8'hEF;
                    16'h94DC: data_out = 8'hF0;
                    16'h94DD: data_out = 8'hF1;
                    16'h94DE: data_out = 8'hF2;
                    16'h94DF: data_out = 8'hF3;
                    16'h94E0: data_out = 8'hF4;
                    16'h94E1: data_out = 8'hF5;
                    16'h94E2: data_out = 8'hF6;
                    16'h94E3: data_out = 8'hF7;
                    16'h94E4: data_out = 8'hF8;
                    16'h94E5: data_out = 8'hF9;
                    16'h94E6: data_out = 8'hFA;
                    16'h94E7: data_out = 8'hFB;
                    16'h94E8: data_out = 8'hFC;
                    16'h94E9: data_out = 8'hFD;
                    16'h94EA: data_out = 8'hFE;
                    16'h94EB: data_out = 8'hFF;
                    16'h94EC: data_out = 8'h80;
                    16'h94ED: data_out = 8'h81;
                    16'h94EE: data_out = 8'h82;
                    16'h94EF: data_out = 8'h83;
                    16'h94F0: data_out = 8'h84;
                    16'h94F1: data_out = 8'h85;
                    16'h94F2: data_out = 8'h86;
                    16'h94F3: data_out = 8'h87;
                    16'h94F4: data_out = 8'h88;
                    16'h94F5: data_out = 8'h89;
                    16'h94F6: data_out = 8'h8A;
                    16'h94F7: data_out = 8'h8B;
                    16'h94F8: data_out = 8'h8C;
                    16'h94F9: data_out = 8'h8D;
                    16'h94FA: data_out = 8'h8E;
                    16'h94FB: data_out = 8'h8F;
                    16'h94FC: data_out = 8'h90;
                    16'h94FD: data_out = 8'h91;
                    16'h94FE: data_out = 8'h92;
                    16'h94FF: data_out = 8'h93;
                    16'h9500: data_out = 8'h95;
                    16'h9501: data_out = 8'h94;
                    16'h9502: data_out = 8'h93;
                    16'h9503: data_out = 8'h92;
                    16'h9504: data_out = 8'h91;
                    16'h9505: data_out = 8'h90;
                    16'h9506: data_out = 8'h8F;
                    16'h9507: data_out = 8'h8E;
                    16'h9508: data_out = 8'h8D;
                    16'h9509: data_out = 8'h8C;
                    16'h950A: data_out = 8'h8B;
                    16'h950B: data_out = 8'h8A;
                    16'h950C: data_out = 8'h89;
                    16'h950D: data_out = 8'h88;
                    16'h950E: data_out = 8'h87;
                    16'h950F: data_out = 8'h86;
                    16'h9510: data_out = 8'h85;
                    16'h9511: data_out = 8'h84;
                    16'h9512: data_out = 8'h83;
                    16'h9513: data_out = 8'h82;
                    16'h9514: data_out = 8'h81;
                    16'h9515: data_out = 8'h0;
                    16'h9516: data_out = 8'h1;
                    16'h9517: data_out = 8'h2;
                    16'h9518: data_out = 8'h3;
                    16'h9519: data_out = 8'h4;
                    16'h951A: data_out = 8'h5;
                    16'h951B: data_out = 8'h6;
                    16'h951C: data_out = 8'h7;
                    16'h951D: data_out = 8'h8;
                    16'h951E: data_out = 8'h9;
                    16'h951F: data_out = 8'hA;
                    16'h9520: data_out = 8'hB;
                    16'h9521: data_out = 8'hC;
                    16'h9522: data_out = 8'hD;
                    16'h9523: data_out = 8'hE;
                    16'h9524: data_out = 8'hF;
                    16'h9525: data_out = 8'h10;
                    16'h9526: data_out = 8'h11;
                    16'h9527: data_out = 8'h12;
                    16'h9528: data_out = 8'h13;
                    16'h9529: data_out = 8'h14;
                    16'h952A: data_out = 8'h15;
                    16'h952B: data_out = 8'h16;
                    16'h952C: data_out = 8'h17;
                    16'h952D: data_out = 8'h18;
                    16'h952E: data_out = 8'h19;
                    16'h952F: data_out = 8'h1A;
                    16'h9530: data_out = 8'h1B;
                    16'h9531: data_out = 8'h1C;
                    16'h9532: data_out = 8'h1D;
                    16'h9533: data_out = 8'h1E;
                    16'h9534: data_out = 8'h1F;
                    16'h9535: data_out = 8'h20;
                    16'h9536: data_out = 8'h21;
                    16'h9537: data_out = 8'h22;
                    16'h9538: data_out = 8'h23;
                    16'h9539: data_out = 8'h24;
                    16'h953A: data_out = 8'h25;
                    16'h953B: data_out = 8'h26;
                    16'h953C: data_out = 8'h27;
                    16'h953D: data_out = 8'h28;
                    16'h953E: data_out = 8'h29;
                    16'h953F: data_out = 8'h2A;
                    16'h9540: data_out = 8'h2B;
                    16'h9541: data_out = 8'h2C;
                    16'h9542: data_out = 8'h2D;
                    16'h9543: data_out = 8'h2E;
                    16'h9544: data_out = 8'h2F;
                    16'h9545: data_out = 8'h30;
                    16'h9546: data_out = 8'h31;
                    16'h9547: data_out = 8'h32;
                    16'h9548: data_out = 8'h33;
                    16'h9549: data_out = 8'h34;
                    16'h954A: data_out = 8'h35;
                    16'h954B: data_out = 8'h36;
                    16'h954C: data_out = 8'h37;
                    16'h954D: data_out = 8'h38;
                    16'h954E: data_out = 8'h39;
                    16'h954F: data_out = 8'h3A;
                    16'h9550: data_out = 8'h3B;
                    16'h9551: data_out = 8'h3C;
                    16'h9552: data_out = 8'h3D;
                    16'h9553: data_out = 8'h3E;
                    16'h9554: data_out = 8'h3F;
                    16'h9555: data_out = 8'h40;
                    16'h9556: data_out = 8'h41;
                    16'h9557: data_out = 8'h42;
                    16'h9558: data_out = 8'h43;
                    16'h9559: data_out = 8'h44;
                    16'h955A: data_out = 8'h45;
                    16'h955B: data_out = 8'h46;
                    16'h955C: data_out = 8'h47;
                    16'h955D: data_out = 8'h48;
                    16'h955E: data_out = 8'h49;
                    16'h955F: data_out = 8'h4A;
                    16'h9560: data_out = 8'h4B;
                    16'h9561: data_out = 8'h4C;
                    16'h9562: data_out = 8'h4D;
                    16'h9563: data_out = 8'h4E;
                    16'h9564: data_out = 8'h4F;
                    16'h9565: data_out = 8'h50;
                    16'h9566: data_out = 8'h51;
                    16'h9567: data_out = 8'h52;
                    16'h9568: data_out = 8'h53;
                    16'h9569: data_out = 8'h54;
                    16'h956A: data_out = 8'h55;
                    16'h956B: data_out = 8'h56;
                    16'h956C: data_out = 8'h57;
                    16'h956D: data_out = 8'h58;
                    16'h956E: data_out = 8'h59;
                    16'h956F: data_out = 8'h5A;
                    16'h9570: data_out = 8'h5B;
                    16'h9571: data_out = 8'h5C;
                    16'h9572: data_out = 8'h5D;
                    16'h9573: data_out = 8'h5E;
                    16'h9574: data_out = 8'h5F;
                    16'h9575: data_out = 8'h60;
                    16'h9576: data_out = 8'h61;
                    16'h9577: data_out = 8'h62;
                    16'h9578: data_out = 8'h63;
                    16'h9579: data_out = 8'h64;
                    16'h957A: data_out = 8'h65;
                    16'h957B: data_out = 8'h66;
                    16'h957C: data_out = 8'h67;
                    16'h957D: data_out = 8'h68;
                    16'h957E: data_out = 8'h69;
                    16'h957F: data_out = 8'h6A;
                    16'h9580: data_out = 8'h95;
                    16'h9581: data_out = 8'h96;
                    16'h9582: data_out = 8'h97;
                    16'h9583: data_out = 8'h98;
                    16'h9584: data_out = 8'h99;
                    16'h9585: data_out = 8'h9A;
                    16'h9586: data_out = 8'h9B;
                    16'h9587: data_out = 8'h9C;
                    16'h9588: data_out = 8'h9D;
                    16'h9589: data_out = 8'h9E;
                    16'h958A: data_out = 8'h9F;
                    16'h958B: data_out = 8'hA0;
                    16'h958C: data_out = 8'hA1;
                    16'h958D: data_out = 8'hA2;
                    16'h958E: data_out = 8'hA3;
                    16'h958F: data_out = 8'hA4;
                    16'h9590: data_out = 8'hA5;
                    16'h9591: data_out = 8'hA6;
                    16'h9592: data_out = 8'hA7;
                    16'h9593: data_out = 8'hA8;
                    16'h9594: data_out = 8'hA9;
                    16'h9595: data_out = 8'hAA;
                    16'h9596: data_out = 8'hAB;
                    16'h9597: data_out = 8'hAC;
                    16'h9598: data_out = 8'hAD;
                    16'h9599: data_out = 8'hAE;
                    16'h959A: data_out = 8'hAF;
                    16'h959B: data_out = 8'hB0;
                    16'h959C: data_out = 8'hB1;
                    16'h959D: data_out = 8'hB2;
                    16'h959E: data_out = 8'hB3;
                    16'h959F: data_out = 8'hB4;
                    16'h95A0: data_out = 8'hB5;
                    16'h95A1: data_out = 8'hB6;
                    16'h95A2: data_out = 8'hB7;
                    16'h95A3: data_out = 8'hB8;
                    16'h95A4: data_out = 8'hB9;
                    16'h95A5: data_out = 8'hBA;
                    16'h95A6: data_out = 8'hBB;
                    16'h95A7: data_out = 8'hBC;
                    16'h95A8: data_out = 8'hBD;
                    16'h95A9: data_out = 8'hBE;
                    16'h95AA: data_out = 8'hBF;
                    16'h95AB: data_out = 8'hC0;
                    16'h95AC: data_out = 8'hC1;
                    16'h95AD: data_out = 8'hC2;
                    16'h95AE: data_out = 8'hC3;
                    16'h95AF: data_out = 8'hC4;
                    16'h95B0: data_out = 8'hC5;
                    16'h95B1: data_out = 8'hC6;
                    16'h95B2: data_out = 8'hC7;
                    16'h95B3: data_out = 8'hC8;
                    16'h95B4: data_out = 8'hC9;
                    16'h95B5: data_out = 8'hCA;
                    16'h95B6: data_out = 8'hCB;
                    16'h95B7: data_out = 8'hCC;
                    16'h95B8: data_out = 8'hCD;
                    16'h95B9: data_out = 8'hCE;
                    16'h95BA: data_out = 8'hCF;
                    16'h95BB: data_out = 8'hD0;
                    16'h95BC: data_out = 8'hD1;
                    16'h95BD: data_out = 8'hD2;
                    16'h95BE: data_out = 8'hD3;
                    16'h95BF: data_out = 8'hD4;
                    16'h95C0: data_out = 8'hD5;
                    16'h95C1: data_out = 8'hD6;
                    16'h95C2: data_out = 8'hD7;
                    16'h95C3: data_out = 8'hD8;
                    16'h95C4: data_out = 8'hD9;
                    16'h95C5: data_out = 8'hDA;
                    16'h95C6: data_out = 8'hDB;
                    16'h95C7: data_out = 8'hDC;
                    16'h95C8: data_out = 8'hDD;
                    16'h95C9: data_out = 8'hDE;
                    16'h95CA: data_out = 8'hDF;
                    16'h95CB: data_out = 8'hE0;
                    16'h95CC: data_out = 8'hE1;
                    16'h95CD: data_out = 8'hE2;
                    16'h95CE: data_out = 8'hE3;
                    16'h95CF: data_out = 8'hE4;
                    16'h95D0: data_out = 8'hE5;
                    16'h95D1: data_out = 8'hE6;
                    16'h95D2: data_out = 8'hE7;
                    16'h95D3: data_out = 8'hE8;
                    16'h95D4: data_out = 8'hE9;
                    16'h95D5: data_out = 8'hEA;
                    16'h95D6: data_out = 8'hEB;
                    16'h95D7: data_out = 8'hEC;
                    16'h95D8: data_out = 8'hED;
                    16'h95D9: data_out = 8'hEE;
                    16'h95DA: data_out = 8'hEF;
                    16'h95DB: data_out = 8'hF0;
                    16'h95DC: data_out = 8'hF1;
                    16'h95DD: data_out = 8'hF2;
                    16'h95DE: data_out = 8'hF3;
                    16'h95DF: data_out = 8'hF4;
                    16'h95E0: data_out = 8'hF5;
                    16'h95E1: data_out = 8'hF6;
                    16'h95E2: data_out = 8'hF7;
                    16'h95E3: data_out = 8'hF8;
                    16'h95E4: data_out = 8'hF9;
                    16'h95E5: data_out = 8'hFA;
                    16'h95E6: data_out = 8'hFB;
                    16'h95E7: data_out = 8'hFC;
                    16'h95E8: data_out = 8'hFD;
                    16'h95E9: data_out = 8'hFE;
                    16'h95EA: data_out = 8'hFF;
                    16'h95EB: data_out = 8'h80;
                    16'h95EC: data_out = 8'h81;
                    16'h95ED: data_out = 8'h82;
                    16'h95EE: data_out = 8'h83;
                    16'h95EF: data_out = 8'h84;
                    16'h95F0: data_out = 8'h85;
                    16'h95F1: data_out = 8'h86;
                    16'h95F2: data_out = 8'h87;
                    16'h95F3: data_out = 8'h88;
                    16'h95F4: data_out = 8'h89;
                    16'h95F5: data_out = 8'h8A;
                    16'h95F6: data_out = 8'h8B;
                    16'h95F7: data_out = 8'h8C;
                    16'h95F8: data_out = 8'h8D;
                    16'h95F9: data_out = 8'h8E;
                    16'h95FA: data_out = 8'h8F;
                    16'h95FB: data_out = 8'h90;
                    16'h95FC: data_out = 8'h91;
                    16'h95FD: data_out = 8'h92;
                    16'h95FE: data_out = 8'h93;
                    16'h95FF: data_out = 8'h94;
                    16'h9600: data_out = 8'h96;
                    16'h9601: data_out = 8'h95;
                    16'h9602: data_out = 8'h94;
                    16'h9603: data_out = 8'h93;
                    16'h9604: data_out = 8'h92;
                    16'h9605: data_out = 8'h91;
                    16'h9606: data_out = 8'h90;
                    16'h9607: data_out = 8'h8F;
                    16'h9608: data_out = 8'h8E;
                    16'h9609: data_out = 8'h8D;
                    16'h960A: data_out = 8'h8C;
                    16'h960B: data_out = 8'h8B;
                    16'h960C: data_out = 8'h8A;
                    16'h960D: data_out = 8'h89;
                    16'h960E: data_out = 8'h88;
                    16'h960F: data_out = 8'h87;
                    16'h9610: data_out = 8'h86;
                    16'h9611: data_out = 8'h85;
                    16'h9612: data_out = 8'h84;
                    16'h9613: data_out = 8'h83;
                    16'h9614: data_out = 8'h82;
                    16'h9615: data_out = 8'h81;
                    16'h9616: data_out = 8'h0;
                    16'h9617: data_out = 8'h1;
                    16'h9618: data_out = 8'h2;
                    16'h9619: data_out = 8'h3;
                    16'h961A: data_out = 8'h4;
                    16'h961B: data_out = 8'h5;
                    16'h961C: data_out = 8'h6;
                    16'h961D: data_out = 8'h7;
                    16'h961E: data_out = 8'h8;
                    16'h961F: data_out = 8'h9;
                    16'h9620: data_out = 8'hA;
                    16'h9621: data_out = 8'hB;
                    16'h9622: data_out = 8'hC;
                    16'h9623: data_out = 8'hD;
                    16'h9624: data_out = 8'hE;
                    16'h9625: data_out = 8'hF;
                    16'h9626: data_out = 8'h10;
                    16'h9627: data_out = 8'h11;
                    16'h9628: data_out = 8'h12;
                    16'h9629: data_out = 8'h13;
                    16'h962A: data_out = 8'h14;
                    16'h962B: data_out = 8'h15;
                    16'h962C: data_out = 8'h16;
                    16'h962D: data_out = 8'h17;
                    16'h962E: data_out = 8'h18;
                    16'h962F: data_out = 8'h19;
                    16'h9630: data_out = 8'h1A;
                    16'h9631: data_out = 8'h1B;
                    16'h9632: data_out = 8'h1C;
                    16'h9633: data_out = 8'h1D;
                    16'h9634: data_out = 8'h1E;
                    16'h9635: data_out = 8'h1F;
                    16'h9636: data_out = 8'h20;
                    16'h9637: data_out = 8'h21;
                    16'h9638: data_out = 8'h22;
                    16'h9639: data_out = 8'h23;
                    16'h963A: data_out = 8'h24;
                    16'h963B: data_out = 8'h25;
                    16'h963C: data_out = 8'h26;
                    16'h963D: data_out = 8'h27;
                    16'h963E: data_out = 8'h28;
                    16'h963F: data_out = 8'h29;
                    16'h9640: data_out = 8'h2A;
                    16'h9641: data_out = 8'h2B;
                    16'h9642: data_out = 8'h2C;
                    16'h9643: data_out = 8'h2D;
                    16'h9644: data_out = 8'h2E;
                    16'h9645: data_out = 8'h2F;
                    16'h9646: data_out = 8'h30;
                    16'h9647: data_out = 8'h31;
                    16'h9648: data_out = 8'h32;
                    16'h9649: data_out = 8'h33;
                    16'h964A: data_out = 8'h34;
                    16'h964B: data_out = 8'h35;
                    16'h964C: data_out = 8'h36;
                    16'h964D: data_out = 8'h37;
                    16'h964E: data_out = 8'h38;
                    16'h964F: data_out = 8'h39;
                    16'h9650: data_out = 8'h3A;
                    16'h9651: data_out = 8'h3B;
                    16'h9652: data_out = 8'h3C;
                    16'h9653: data_out = 8'h3D;
                    16'h9654: data_out = 8'h3E;
                    16'h9655: data_out = 8'h3F;
                    16'h9656: data_out = 8'h40;
                    16'h9657: data_out = 8'h41;
                    16'h9658: data_out = 8'h42;
                    16'h9659: data_out = 8'h43;
                    16'h965A: data_out = 8'h44;
                    16'h965B: data_out = 8'h45;
                    16'h965C: data_out = 8'h46;
                    16'h965D: data_out = 8'h47;
                    16'h965E: data_out = 8'h48;
                    16'h965F: data_out = 8'h49;
                    16'h9660: data_out = 8'h4A;
                    16'h9661: data_out = 8'h4B;
                    16'h9662: data_out = 8'h4C;
                    16'h9663: data_out = 8'h4D;
                    16'h9664: data_out = 8'h4E;
                    16'h9665: data_out = 8'h4F;
                    16'h9666: data_out = 8'h50;
                    16'h9667: data_out = 8'h51;
                    16'h9668: data_out = 8'h52;
                    16'h9669: data_out = 8'h53;
                    16'h966A: data_out = 8'h54;
                    16'h966B: data_out = 8'h55;
                    16'h966C: data_out = 8'h56;
                    16'h966D: data_out = 8'h57;
                    16'h966E: data_out = 8'h58;
                    16'h966F: data_out = 8'h59;
                    16'h9670: data_out = 8'h5A;
                    16'h9671: data_out = 8'h5B;
                    16'h9672: data_out = 8'h5C;
                    16'h9673: data_out = 8'h5D;
                    16'h9674: data_out = 8'h5E;
                    16'h9675: data_out = 8'h5F;
                    16'h9676: data_out = 8'h60;
                    16'h9677: data_out = 8'h61;
                    16'h9678: data_out = 8'h62;
                    16'h9679: data_out = 8'h63;
                    16'h967A: data_out = 8'h64;
                    16'h967B: data_out = 8'h65;
                    16'h967C: data_out = 8'h66;
                    16'h967D: data_out = 8'h67;
                    16'h967E: data_out = 8'h68;
                    16'h967F: data_out = 8'h69;
                    16'h9680: data_out = 8'h96;
                    16'h9681: data_out = 8'h97;
                    16'h9682: data_out = 8'h98;
                    16'h9683: data_out = 8'h99;
                    16'h9684: data_out = 8'h9A;
                    16'h9685: data_out = 8'h9B;
                    16'h9686: data_out = 8'h9C;
                    16'h9687: data_out = 8'h9D;
                    16'h9688: data_out = 8'h9E;
                    16'h9689: data_out = 8'h9F;
                    16'h968A: data_out = 8'hA0;
                    16'h968B: data_out = 8'hA1;
                    16'h968C: data_out = 8'hA2;
                    16'h968D: data_out = 8'hA3;
                    16'h968E: data_out = 8'hA4;
                    16'h968F: data_out = 8'hA5;
                    16'h9690: data_out = 8'hA6;
                    16'h9691: data_out = 8'hA7;
                    16'h9692: data_out = 8'hA8;
                    16'h9693: data_out = 8'hA9;
                    16'h9694: data_out = 8'hAA;
                    16'h9695: data_out = 8'hAB;
                    16'h9696: data_out = 8'hAC;
                    16'h9697: data_out = 8'hAD;
                    16'h9698: data_out = 8'hAE;
                    16'h9699: data_out = 8'hAF;
                    16'h969A: data_out = 8'hB0;
                    16'h969B: data_out = 8'hB1;
                    16'h969C: data_out = 8'hB2;
                    16'h969D: data_out = 8'hB3;
                    16'h969E: data_out = 8'hB4;
                    16'h969F: data_out = 8'hB5;
                    16'h96A0: data_out = 8'hB6;
                    16'h96A1: data_out = 8'hB7;
                    16'h96A2: data_out = 8'hB8;
                    16'h96A3: data_out = 8'hB9;
                    16'h96A4: data_out = 8'hBA;
                    16'h96A5: data_out = 8'hBB;
                    16'h96A6: data_out = 8'hBC;
                    16'h96A7: data_out = 8'hBD;
                    16'h96A8: data_out = 8'hBE;
                    16'h96A9: data_out = 8'hBF;
                    16'h96AA: data_out = 8'hC0;
                    16'h96AB: data_out = 8'hC1;
                    16'h96AC: data_out = 8'hC2;
                    16'h96AD: data_out = 8'hC3;
                    16'h96AE: data_out = 8'hC4;
                    16'h96AF: data_out = 8'hC5;
                    16'h96B0: data_out = 8'hC6;
                    16'h96B1: data_out = 8'hC7;
                    16'h96B2: data_out = 8'hC8;
                    16'h96B3: data_out = 8'hC9;
                    16'h96B4: data_out = 8'hCA;
                    16'h96B5: data_out = 8'hCB;
                    16'h96B6: data_out = 8'hCC;
                    16'h96B7: data_out = 8'hCD;
                    16'h96B8: data_out = 8'hCE;
                    16'h96B9: data_out = 8'hCF;
                    16'h96BA: data_out = 8'hD0;
                    16'h96BB: data_out = 8'hD1;
                    16'h96BC: data_out = 8'hD2;
                    16'h96BD: data_out = 8'hD3;
                    16'h96BE: data_out = 8'hD4;
                    16'h96BF: data_out = 8'hD5;
                    16'h96C0: data_out = 8'hD6;
                    16'h96C1: data_out = 8'hD7;
                    16'h96C2: data_out = 8'hD8;
                    16'h96C3: data_out = 8'hD9;
                    16'h96C4: data_out = 8'hDA;
                    16'h96C5: data_out = 8'hDB;
                    16'h96C6: data_out = 8'hDC;
                    16'h96C7: data_out = 8'hDD;
                    16'h96C8: data_out = 8'hDE;
                    16'h96C9: data_out = 8'hDF;
                    16'h96CA: data_out = 8'hE0;
                    16'h96CB: data_out = 8'hE1;
                    16'h96CC: data_out = 8'hE2;
                    16'h96CD: data_out = 8'hE3;
                    16'h96CE: data_out = 8'hE4;
                    16'h96CF: data_out = 8'hE5;
                    16'h96D0: data_out = 8'hE6;
                    16'h96D1: data_out = 8'hE7;
                    16'h96D2: data_out = 8'hE8;
                    16'h96D3: data_out = 8'hE9;
                    16'h96D4: data_out = 8'hEA;
                    16'h96D5: data_out = 8'hEB;
                    16'h96D6: data_out = 8'hEC;
                    16'h96D7: data_out = 8'hED;
                    16'h96D8: data_out = 8'hEE;
                    16'h96D9: data_out = 8'hEF;
                    16'h96DA: data_out = 8'hF0;
                    16'h96DB: data_out = 8'hF1;
                    16'h96DC: data_out = 8'hF2;
                    16'h96DD: data_out = 8'hF3;
                    16'h96DE: data_out = 8'hF4;
                    16'h96DF: data_out = 8'hF5;
                    16'h96E0: data_out = 8'hF6;
                    16'h96E1: data_out = 8'hF7;
                    16'h96E2: data_out = 8'hF8;
                    16'h96E3: data_out = 8'hF9;
                    16'h96E4: data_out = 8'hFA;
                    16'h96E5: data_out = 8'hFB;
                    16'h96E6: data_out = 8'hFC;
                    16'h96E7: data_out = 8'hFD;
                    16'h96E8: data_out = 8'hFE;
                    16'h96E9: data_out = 8'hFF;
                    16'h96EA: data_out = 8'h80;
                    16'h96EB: data_out = 8'h81;
                    16'h96EC: data_out = 8'h82;
                    16'h96ED: data_out = 8'h83;
                    16'h96EE: data_out = 8'h84;
                    16'h96EF: data_out = 8'h85;
                    16'h96F0: data_out = 8'h86;
                    16'h96F1: data_out = 8'h87;
                    16'h96F2: data_out = 8'h88;
                    16'h96F3: data_out = 8'h89;
                    16'h96F4: data_out = 8'h8A;
                    16'h96F5: data_out = 8'h8B;
                    16'h96F6: data_out = 8'h8C;
                    16'h96F7: data_out = 8'h8D;
                    16'h96F8: data_out = 8'h8E;
                    16'h96F9: data_out = 8'h8F;
                    16'h96FA: data_out = 8'h90;
                    16'h96FB: data_out = 8'h91;
                    16'h96FC: data_out = 8'h92;
                    16'h96FD: data_out = 8'h93;
                    16'h96FE: data_out = 8'h94;
                    16'h96FF: data_out = 8'h95;
                    16'h9700: data_out = 8'h97;
                    16'h9701: data_out = 8'h96;
                    16'h9702: data_out = 8'h95;
                    16'h9703: data_out = 8'h94;
                    16'h9704: data_out = 8'h93;
                    16'h9705: data_out = 8'h92;
                    16'h9706: data_out = 8'h91;
                    16'h9707: data_out = 8'h90;
                    16'h9708: data_out = 8'h8F;
                    16'h9709: data_out = 8'h8E;
                    16'h970A: data_out = 8'h8D;
                    16'h970B: data_out = 8'h8C;
                    16'h970C: data_out = 8'h8B;
                    16'h970D: data_out = 8'h8A;
                    16'h970E: data_out = 8'h89;
                    16'h970F: data_out = 8'h88;
                    16'h9710: data_out = 8'h87;
                    16'h9711: data_out = 8'h86;
                    16'h9712: data_out = 8'h85;
                    16'h9713: data_out = 8'h84;
                    16'h9714: data_out = 8'h83;
                    16'h9715: data_out = 8'h82;
                    16'h9716: data_out = 8'h81;
                    16'h9717: data_out = 8'h0;
                    16'h9718: data_out = 8'h1;
                    16'h9719: data_out = 8'h2;
                    16'h971A: data_out = 8'h3;
                    16'h971B: data_out = 8'h4;
                    16'h971C: data_out = 8'h5;
                    16'h971D: data_out = 8'h6;
                    16'h971E: data_out = 8'h7;
                    16'h971F: data_out = 8'h8;
                    16'h9720: data_out = 8'h9;
                    16'h9721: data_out = 8'hA;
                    16'h9722: data_out = 8'hB;
                    16'h9723: data_out = 8'hC;
                    16'h9724: data_out = 8'hD;
                    16'h9725: data_out = 8'hE;
                    16'h9726: data_out = 8'hF;
                    16'h9727: data_out = 8'h10;
                    16'h9728: data_out = 8'h11;
                    16'h9729: data_out = 8'h12;
                    16'h972A: data_out = 8'h13;
                    16'h972B: data_out = 8'h14;
                    16'h972C: data_out = 8'h15;
                    16'h972D: data_out = 8'h16;
                    16'h972E: data_out = 8'h17;
                    16'h972F: data_out = 8'h18;
                    16'h9730: data_out = 8'h19;
                    16'h9731: data_out = 8'h1A;
                    16'h9732: data_out = 8'h1B;
                    16'h9733: data_out = 8'h1C;
                    16'h9734: data_out = 8'h1D;
                    16'h9735: data_out = 8'h1E;
                    16'h9736: data_out = 8'h1F;
                    16'h9737: data_out = 8'h20;
                    16'h9738: data_out = 8'h21;
                    16'h9739: data_out = 8'h22;
                    16'h973A: data_out = 8'h23;
                    16'h973B: data_out = 8'h24;
                    16'h973C: data_out = 8'h25;
                    16'h973D: data_out = 8'h26;
                    16'h973E: data_out = 8'h27;
                    16'h973F: data_out = 8'h28;
                    16'h9740: data_out = 8'h29;
                    16'h9741: data_out = 8'h2A;
                    16'h9742: data_out = 8'h2B;
                    16'h9743: data_out = 8'h2C;
                    16'h9744: data_out = 8'h2D;
                    16'h9745: data_out = 8'h2E;
                    16'h9746: data_out = 8'h2F;
                    16'h9747: data_out = 8'h30;
                    16'h9748: data_out = 8'h31;
                    16'h9749: data_out = 8'h32;
                    16'h974A: data_out = 8'h33;
                    16'h974B: data_out = 8'h34;
                    16'h974C: data_out = 8'h35;
                    16'h974D: data_out = 8'h36;
                    16'h974E: data_out = 8'h37;
                    16'h974F: data_out = 8'h38;
                    16'h9750: data_out = 8'h39;
                    16'h9751: data_out = 8'h3A;
                    16'h9752: data_out = 8'h3B;
                    16'h9753: data_out = 8'h3C;
                    16'h9754: data_out = 8'h3D;
                    16'h9755: data_out = 8'h3E;
                    16'h9756: data_out = 8'h3F;
                    16'h9757: data_out = 8'h40;
                    16'h9758: data_out = 8'h41;
                    16'h9759: data_out = 8'h42;
                    16'h975A: data_out = 8'h43;
                    16'h975B: data_out = 8'h44;
                    16'h975C: data_out = 8'h45;
                    16'h975D: data_out = 8'h46;
                    16'h975E: data_out = 8'h47;
                    16'h975F: data_out = 8'h48;
                    16'h9760: data_out = 8'h49;
                    16'h9761: data_out = 8'h4A;
                    16'h9762: data_out = 8'h4B;
                    16'h9763: data_out = 8'h4C;
                    16'h9764: data_out = 8'h4D;
                    16'h9765: data_out = 8'h4E;
                    16'h9766: data_out = 8'h4F;
                    16'h9767: data_out = 8'h50;
                    16'h9768: data_out = 8'h51;
                    16'h9769: data_out = 8'h52;
                    16'h976A: data_out = 8'h53;
                    16'h976B: data_out = 8'h54;
                    16'h976C: data_out = 8'h55;
                    16'h976D: data_out = 8'h56;
                    16'h976E: data_out = 8'h57;
                    16'h976F: data_out = 8'h58;
                    16'h9770: data_out = 8'h59;
                    16'h9771: data_out = 8'h5A;
                    16'h9772: data_out = 8'h5B;
                    16'h9773: data_out = 8'h5C;
                    16'h9774: data_out = 8'h5D;
                    16'h9775: data_out = 8'h5E;
                    16'h9776: data_out = 8'h5F;
                    16'h9777: data_out = 8'h60;
                    16'h9778: data_out = 8'h61;
                    16'h9779: data_out = 8'h62;
                    16'h977A: data_out = 8'h63;
                    16'h977B: data_out = 8'h64;
                    16'h977C: data_out = 8'h65;
                    16'h977D: data_out = 8'h66;
                    16'h977E: data_out = 8'h67;
                    16'h977F: data_out = 8'h68;
                    16'h9780: data_out = 8'h97;
                    16'h9781: data_out = 8'h98;
                    16'h9782: data_out = 8'h99;
                    16'h9783: data_out = 8'h9A;
                    16'h9784: data_out = 8'h9B;
                    16'h9785: data_out = 8'h9C;
                    16'h9786: data_out = 8'h9D;
                    16'h9787: data_out = 8'h9E;
                    16'h9788: data_out = 8'h9F;
                    16'h9789: data_out = 8'hA0;
                    16'h978A: data_out = 8'hA1;
                    16'h978B: data_out = 8'hA2;
                    16'h978C: data_out = 8'hA3;
                    16'h978D: data_out = 8'hA4;
                    16'h978E: data_out = 8'hA5;
                    16'h978F: data_out = 8'hA6;
                    16'h9790: data_out = 8'hA7;
                    16'h9791: data_out = 8'hA8;
                    16'h9792: data_out = 8'hA9;
                    16'h9793: data_out = 8'hAA;
                    16'h9794: data_out = 8'hAB;
                    16'h9795: data_out = 8'hAC;
                    16'h9796: data_out = 8'hAD;
                    16'h9797: data_out = 8'hAE;
                    16'h9798: data_out = 8'hAF;
                    16'h9799: data_out = 8'hB0;
                    16'h979A: data_out = 8'hB1;
                    16'h979B: data_out = 8'hB2;
                    16'h979C: data_out = 8'hB3;
                    16'h979D: data_out = 8'hB4;
                    16'h979E: data_out = 8'hB5;
                    16'h979F: data_out = 8'hB6;
                    16'h97A0: data_out = 8'hB7;
                    16'h97A1: data_out = 8'hB8;
                    16'h97A2: data_out = 8'hB9;
                    16'h97A3: data_out = 8'hBA;
                    16'h97A4: data_out = 8'hBB;
                    16'h97A5: data_out = 8'hBC;
                    16'h97A6: data_out = 8'hBD;
                    16'h97A7: data_out = 8'hBE;
                    16'h97A8: data_out = 8'hBF;
                    16'h97A9: data_out = 8'hC0;
                    16'h97AA: data_out = 8'hC1;
                    16'h97AB: data_out = 8'hC2;
                    16'h97AC: data_out = 8'hC3;
                    16'h97AD: data_out = 8'hC4;
                    16'h97AE: data_out = 8'hC5;
                    16'h97AF: data_out = 8'hC6;
                    16'h97B0: data_out = 8'hC7;
                    16'h97B1: data_out = 8'hC8;
                    16'h97B2: data_out = 8'hC9;
                    16'h97B3: data_out = 8'hCA;
                    16'h97B4: data_out = 8'hCB;
                    16'h97B5: data_out = 8'hCC;
                    16'h97B6: data_out = 8'hCD;
                    16'h97B7: data_out = 8'hCE;
                    16'h97B8: data_out = 8'hCF;
                    16'h97B9: data_out = 8'hD0;
                    16'h97BA: data_out = 8'hD1;
                    16'h97BB: data_out = 8'hD2;
                    16'h97BC: data_out = 8'hD3;
                    16'h97BD: data_out = 8'hD4;
                    16'h97BE: data_out = 8'hD5;
                    16'h97BF: data_out = 8'hD6;
                    16'h97C0: data_out = 8'hD7;
                    16'h97C1: data_out = 8'hD8;
                    16'h97C2: data_out = 8'hD9;
                    16'h97C3: data_out = 8'hDA;
                    16'h97C4: data_out = 8'hDB;
                    16'h97C5: data_out = 8'hDC;
                    16'h97C6: data_out = 8'hDD;
                    16'h97C7: data_out = 8'hDE;
                    16'h97C8: data_out = 8'hDF;
                    16'h97C9: data_out = 8'hE0;
                    16'h97CA: data_out = 8'hE1;
                    16'h97CB: data_out = 8'hE2;
                    16'h97CC: data_out = 8'hE3;
                    16'h97CD: data_out = 8'hE4;
                    16'h97CE: data_out = 8'hE5;
                    16'h97CF: data_out = 8'hE6;
                    16'h97D0: data_out = 8'hE7;
                    16'h97D1: data_out = 8'hE8;
                    16'h97D2: data_out = 8'hE9;
                    16'h97D3: data_out = 8'hEA;
                    16'h97D4: data_out = 8'hEB;
                    16'h97D5: data_out = 8'hEC;
                    16'h97D6: data_out = 8'hED;
                    16'h97D7: data_out = 8'hEE;
                    16'h97D8: data_out = 8'hEF;
                    16'h97D9: data_out = 8'hF0;
                    16'h97DA: data_out = 8'hF1;
                    16'h97DB: data_out = 8'hF2;
                    16'h97DC: data_out = 8'hF3;
                    16'h97DD: data_out = 8'hF4;
                    16'h97DE: data_out = 8'hF5;
                    16'h97DF: data_out = 8'hF6;
                    16'h97E0: data_out = 8'hF7;
                    16'h97E1: data_out = 8'hF8;
                    16'h97E2: data_out = 8'hF9;
                    16'h97E3: data_out = 8'hFA;
                    16'h97E4: data_out = 8'hFB;
                    16'h97E5: data_out = 8'hFC;
                    16'h97E6: data_out = 8'hFD;
                    16'h97E7: data_out = 8'hFE;
                    16'h97E8: data_out = 8'hFF;
                    16'h97E9: data_out = 8'h80;
                    16'h97EA: data_out = 8'h81;
                    16'h97EB: data_out = 8'h82;
                    16'h97EC: data_out = 8'h83;
                    16'h97ED: data_out = 8'h84;
                    16'h97EE: data_out = 8'h85;
                    16'h97EF: data_out = 8'h86;
                    16'h97F0: data_out = 8'h87;
                    16'h97F1: data_out = 8'h88;
                    16'h97F2: data_out = 8'h89;
                    16'h97F3: data_out = 8'h8A;
                    16'h97F4: data_out = 8'h8B;
                    16'h97F5: data_out = 8'h8C;
                    16'h97F6: data_out = 8'h8D;
                    16'h97F7: data_out = 8'h8E;
                    16'h97F8: data_out = 8'h8F;
                    16'h97F9: data_out = 8'h90;
                    16'h97FA: data_out = 8'h91;
                    16'h97FB: data_out = 8'h92;
                    16'h97FC: data_out = 8'h93;
                    16'h97FD: data_out = 8'h94;
                    16'h97FE: data_out = 8'h95;
                    16'h97FF: data_out = 8'h96;
                    16'h9800: data_out = 8'h98;
                    16'h9801: data_out = 8'h97;
                    16'h9802: data_out = 8'h96;
                    16'h9803: data_out = 8'h95;
                    16'h9804: data_out = 8'h94;
                    16'h9805: data_out = 8'h93;
                    16'h9806: data_out = 8'h92;
                    16'h9807: data_out = 8'h91;
                    16'h9808: data_out = 8'h90;
                    16'h9809: data_out = 8'h8F;
                    16'h980A: data_out = 8'h8E;
                    16'h980B: data_out = 8'h8D;
                    16'h980C: data_out = 8'h8C;
                    16'h980D: data_out = 8'h8B;
                    16'h980E: data_out = 8'h8A;
                    16'h980F: data_out = 8'h89;
                    16'h9810: data_out = 8'h88;
                    16'h9811: data_out = 8'h87;
                    16'h9812: data_out = 8'h86;
                    16'h9813: data_out = 8'h85;
                    16'h9814: data_out = 8'h84;
                    16'h9815: data_out = 8'h83;
                    16'h9816: data_out = 8'h82;
                    16'h9817: data_out = 8'h81;
                    16'h9818: data_out = 8'h0;
                    16'h9819: data_out = 8'h1;
                    16'h981A: data_out = 8'h2;
                    16'h981B: data_out = 8'h3;
                    16'h981C: data_out = 8'h4;
                    16'h981D: data_out = 8'h5;
                    16'h981E: data_out = 8'h6;
                    16'h981F: data_out = 8'h7;
                    16'h9820: data_out = 8'h8;
                    16'h9821: data_out = 8'h9;
                    16'h9822: data_out = 8'hA;
                    16'h9823: data_out = 8'hB;
                    16'h9824: data_out = 8'hC;
                    16'h9825: data_out = 8'hD;
                    16'h9826: data_out = 8'hE;
                    16'h9827: data_out = 8'hF;
                    16'h9828: data_out = 8'h10;
                    16'h9829: data_out = 8'h11;
                    16'h982A: data_out = 8'h12;
                    16'h982B: data_out = 8'h13;
                    16'h982C: data_out = 8'h14;
                    16'h982D: data_out = 8'h15;
                    16'h982E: data_out = 8'h16;
                    16'h982F: data_out = 8'h17;
                    16'h9830: data_out = 8'h18;
                    16'h9831: data_out = 8'h19;
                    16'h9832: data_out = 8'h1A;
                    16'h9833: data_out = 8'h1B;
                    16'h9834: data_out = 8'h1C;
                    16'h9835: data_out = 8'h1D;
                    16'h9836: data_out = 8'h1E;
                    16'h9837: data_out = 8'h1F;
                    16'h9838: data_out = 8'h20;
                    16'h9839: data_out = 8'h21;
                    16'h983A: data_out = 8'h22;
                    16'h983B: data_out = 8'h23;
                    16'h983C: data_out = 8'h24;
                    16'h983D: data_out = 8'h25;
                    16'h983E: data_out = 8'h26;
                    16'h983F: data_out = 8'h27;
                    16'h9840: data_out = 8'h28;
                    16'h9841: data_out = 8'h29;
                    16'h9842: data_out = 8'h2A;
                    16'h9843: data_out = 8'h2B;
                    16'h9844: data_out = 8'h2C;
                    16'h9845: data_out = 8'h2D;
                    16'h9846: data_out = 8'h2E;
                    16'h9847: data_out = 8'h2F;
                    16'h9848: data_out = 8'h30;
                    16'h9849: data_out = 8'h31;
                    16'h984A: data_out = 8'h32;
                    16'h984B: data_out = 8'h33;
                    16'h984C: data_out = 8'h34;
                    16'h984D: data_out = 8'h35;
                    16'h984E: data_out = 8'h36;
                    16'h984F: data_out = 8'h37;
                    16'h9850: data_out = 8'h38;
                    16'h9851: data_out = 8'h39;
                    16'h9852: data_out = 8'h3A;
                    16'h9853: data_out = 8'h3B;
                    16'h9854: data_out = 8'h3C;
                    16'h9855: data_out = 8'h3D;
                    16'h9856: data_out = 8'h3E;
                    16'h9857: data_out = 8'h3F;
                    16'h9858: data_out = 8'h40;
                    16'h9859: data_out = 8'h41;
                    16'h985A: data_out = 8'h42;
                    16'h985B: data_out = 8'h43;
                    16'h985C: data_out = 8'h44;
                    16'h985D: data_out = 8'h45;
                    16'h985E: data_out = 8'h46;
                    16'h985F: data_out = 8'h47;
                    16'h9860: data_out = 8'h48;
                    16'h9861: data_out = 8'h49;
                    16'h9862: data_out = 8'h4A;
                    16'h9863: data_out = 8'h4B;
                    16'h9864: data_out = 8'h4C;
                    16'h9865: data_out = 8'h4D;
                    16'h9866: data_out = 8'h4E;
                    16'h9867: data_out = 8'h4F;
                    16'h9868: data_out = 8'h50;
                    16'h9869: data_out = 8'h51;
                    16'h986A: data_out = 8'h52;
                    16'h986B: data_out = 8'h53;
                    16'h986C: data_out = 8'h54;
                    16'h986D: data_out = 8'h55;
                    16'h986E: data_out = 8'h56;
                    16'h986F: data_out = 8'h57;
                    16'h9870: data_out = 8'h58;
                    16'h9871: data_out = 8'h59;
                    16'h9872: data_out = 8'h5A;
                    16'h9873: data_out = 8'h5B;
                    16'h9874: data_out = 8'h5C;
                    16'h9875: data_out = 8'h5D;
                    16'h9876: data_out = 8'h5E;
                    16'h9877: data_out = 8'h5F;
                    16'h9878: data_out = 8'h60;
                    16'h9879: data_out = 8'h61;
                    16'h987A: data_out = 8'h62;
                    16'h987B: data_out = 8'h63;
                    16'h987C: data_out = 8'h64;
                    16'h987D: data_out = 8'h65;
                    16'h987E: data_out = 8'h66;
                    16'h987F: data_out = 8'h67;
                    16'h9880: data_out = 8'h98;
                    16'h9881: data_out = 8'h99;
                    16'h9882: data_out = 8'h9A;
                    16'h9883: data_out = 8'h9B;
                    16'h9884: data_out = 8'h9C;
                    16'h9885: data_out = 8'h9D;
                    16'h9886: data_out = 8'h9E;
                    16'h9887: data_out = 8'h9F;
                    16'h9888: data_out = 8'hA0;
                    16'h9889: data_out = 8'hA1;
                    16'h988A: data_out = 8'hA2;
                    16'h988B: data_out = 8'hA3;
                    16'h988C: data_out = 8'hA4;
                    16'h988D: data_out = 8'hA5;
                    16'h988E: data_out = 8'hA6;
                    16'h988F: data_out = 8'hA7;
                    16'h9890: data_out = 8'hA8;
                    16'h9891: data_out = 8'hA9;
                    16'h9892: data_out = 8'hAA;
                    16'h9893: data_out = 8'hAB;
                    16'h9894: data_out = 8'hAC;
                    16'h9895: data_out = 8'hAD;
                    16'h9896: data_out = 8'hAE;
                    16'h9897: data_out = 8'hAF;
                    16'h9898: data_out = 8'hB0;
                    16'h9899: data_out = 8'hB1;
                    16'h989A: data_out = 8'hB2;
                    16'h989B: data_out = 8'hB3;
                    16'h989C: data_out = 8'hB4;
                    16'h989D: data_out = 8'hB5;
                    16'h989E: data_out = 8'hB6;
                    16'h989F: data_out = 8'hB7;
                    16'h98A0: data_out = 8'hB8;
                    16'h98A1: data_out = 8'hB9;
                    16'h98A2: data_out = 8'hBA;
                    16'h98A3: data_out = 8'hBB;
                    16'h98A4: data_out = 8'hBC;
                    16'h98A5: data_out = 8'hBD;
                    16'h98A6: data_out = 8'hBE;
                    16'h98A7: data_out = 8'hBF;
                    16'h98A8: data_out = 8'hC0;
                    16'h98A9: data_out = 8'hC1;
                    16'h98AA: data_out = 8'hC2;
                    16'h98AB: data_out = 8'hC3;
                    16'h98AC: data_out = 8'hC4;
                    16'h98AD: data_out = 8'hC5;
                    16'h98AE: data_out = 8'hC6;
                    16'h98AF: data_out = 8'hC7;
                    16'h98B0: data_out = 8'hC8;
                    16'h98B1: data_out = 8'hC9;
                    16'h98B2: data_out = 8'hCA;
                    16'h98B3: data_out = 8'hCB;
                    16'h98B4: data_out = 8'hCC;
                    16'h98B5: data_out = 8'hCD;
                    16'h98B6: data_out = 8'hCE;
                    16'h98B7: data_out = 8'hCF;
                    16'h98B8: data_out = 8'hD0;
                    16'h98B9: data_out = 8'hD1;
                    16'h98BA: data_out = 8'hD2;
                    16'h98BB: data_out = 8'hD3;
                    16'h98BC: data_out = 8'hD4;
                    16'h98BD: data_out = 8'hD5;
                    16'h98BE: data_out = 8'hD6;
                    16'h98BF: data_out = 8'hD7;
                    16'h98C0: data_out = 8'hD8;
                    16'h98C1: data_out = 8'hD9;
                    16'h98C2: data_out = 8'hDA;
                    16'h98C3: data_out = 8'hDB;
                    16'h98C4: data_out = 8'hDC;
                    16'h98C5: data_out = 8'hDD;
                    16'h98C6: data_out = 8'hDE;
                    16'h98C7: data_out = 8'hDF;
                    16'h98C8: data_out = 8'hE0;
                    16'h98C9: data_out = 8'hE1;
                    16'h98CA: data_out = 8'hE2;
                    16'h98CB: data_out = 8'hE3;
                    16'h98CC: data_out = 8'hE4;
                    16'h98CD: data_out = 8'hE5;
                    16'h98CE: data_out = 8'hE6;
                    16'h98CF: data_out = 8'hE7;
                    16'h98D0: data_out = 8'hE8;
                    16'h98D1: data_out = 8'hE9;
                    16'h98D2: data_out = 8'hEA;
                    16'h98D3: data_out = 8'hEB;
                    16'h98D4: data_out = 8'hEC;
                    16'h98D5: data_out = 8'hED;
                    16'h98D6: data_out = 8'hEE;
                    16'h98D7: data_out = 8'hEF;
                    16'h98D8: data_out = 8'hF0;
                    16'h98D9: data_out = 8'hF1;
                    16'h98DA: data_out = 8'hF2;
                    16'h98DB: data_out = 8'hF3;
                    16'h98DC: data_out = 8'hF4;
                    16'h98DD: data_out = 8'hF5;
                    16'h98DE: data_out = 8'hF6;
                    16'h98DF: data_out = 8'hF7;
                    16'h98E0: data_out = 8'hF8;
                    16'h98E1: data_out = 8'hF9;
                    16'h98E2: data_out = 8'hFA;
                    16'h98E3: data_out = 8'hFB;
                    16'h98E4: data_out = 8'hFC;
                    16'h98E5: data_out = 8'hFD;
                    16'h98E6: data_out = 8'hFE;
                    16'h98E7: data_out = 8'hFF;
                    16'h98E8: data_out = 8'h80;
                    16'h98E9: data_out = 8'h81;
                    16'h98EA: data_out = 8'h82;
                    16'h98EB: data_out = 8'h83;
                    16'h98EC: data_out = 8'h84;
                    16'h98ED: data_out = 8'h85;
                    16'h98EE: data_out = 8'h86;
                    16'h98EF: data_out = 8'h87;
                    16'h98F0: data_out = 8'h88;
                    16'h98F1: data_out = 8'h89;
                    16'h98F2: data_out = 8'h8A;
                    16'h98F3: data_out = 8'h8B;
                    16'h98F4: data_out = 8'h8C;
                    16'h98F5: data_out = 8'h8D;
                    16'h98F6: data_out = 8'h8E;
                    16'h98F7: data_out = 8'h8F;
                    16'h98F8: data_out = 8'h90;
                    16'h98F9: data_out = 8'h91;
                    16'h98FA: data_out = 8'h92;
                    16'h98FB: data_out = 8'h93;
                    16'h98FC: data_out = 8'h94;
                    16'h98FD: data_out = 8'h95;
                    16'h98FE: data_out = 8'h96;
                    16'h98FF: data_out = 8'h97;
                    16'h9900: data_out = 8'h99;
                    16'h9901: data_out = 8'h98;
                    16'h9902: data_out = 8'h97;
                    16'h9903: data_out = 8'h96;
                    16'h9904: data_out = 8'h95;
                    16'h9905: data_out = 8'h94;
                    16'h9906: data_out = 8'h93;
                    16'h9907: data_out = 8'h92;
                    16'h9908: data_out = 8'h91;
                    16'h9909: data_out = 8'h90;
                    16'h990A: data_out = 8'h8F;
                    16'h990B: data_out = 8'h8E;
                    16'h990C: data_out = 8'h8D;
                    16'h990D: data_out = 8'h8C;
                    16'h990E: data_out = 8'h8B;
                    16'h990F: data_out = 8'h8A;
                    16'h9910: data_out = 8'h89;
                    16'h9911: data_out = 8'h88;
                    16'h9912: data_out = 8'h87;
                    16'h9913: data_out = 8'h86;
                    16'h9914: data_out = 8'h85;
                    16'h9915: data_out = 8'h84;
                    16'h9916: data_out = 8'h83;
                    16'h9917: data_out = 8'h82;
                    16'h9918: data_out = 8'h81;
                    16'h9919: data_out = 8'h0;
                    16'h991A: data_out = 8'h1;
                    16'h991B: data_out = 8'h2;
                    16'h991C: data_out = 8'h3;
                    16'h991D: data_out = 8'h4;
                    16'h991E: data_out = 8'h5;
                    16'h991F: data_out = 8'h6;
                    16'h9920: data_out = 8'h7;
                    16'h9921: data_out = 8'h8;
                    16'h9922: data_out = 8'h9;
                    16'h9923: data_out = 8'hA;
                    16'h9924: data_out = 8'hB;
                    16'h9925: data_out = 8'hC;
                    16'h9926: data_out = 8'hD;
                    16'h9927: data_out = 8'hE;
                    16'h9928: data_out = 8'hF;
                    16'h9929: data_out = 8'h10;
                    16'h992A: data_out = 8'h11;
                    16'h992B: data_out = 8'h12;
                    16'h992C: data_out = 8'h13;
                    16'h992D: data_out = 8'h14;
                    16'h992E: data_out = 8'h15;
                    16'h992F: data_out = 8'h16;
                    16'h9930: data_out = 8'h17;
                    16'h9931: data_out = 8'h18;
                    16'h9932: data_out = 8'h19;
                    16'h9933: data_out = 8'h1A;
                    16'h9934: data_out = 8'h1B;
                    16'h9935: data_out = 8'h1C;
                    16'h9936: data_out = 8'h1D;
                    16'h9937: data_out = 8'h1E;
                    16'h9938: data_out = 8'h1F;
                    16'h9939: data_out = 8'h20;
                    16'h993A: data_out = 8'h21;
                    16'h993B: data_out = 8'h22;
                    16'h993C: data_out = 8'h23;
                    16'h993D: data_out = 8'h24;
                    16'h993E: data_out = 8'h25;
                    16'h993F: data_out = 8'h26;
                    16'h9940: data_out = 8'h27;
                    16'h9941: data_out = 8'h28;
                    16'h9942: data_out = 8'h29;
                    16'h9943: data_out = 8'h2A;
                    16'h9944: data_out = 8'h2B;
                    16'h9945: data_out = 8'h2C;
                    16'h9946: data_out = 8'h2D;
                    16'h9947: data_out = 8'h2E;
                    16'h9948: data_out = 8'h2F;
                    16'h9949: data_out = 8'h30;
                    16'h994A: data_out = 8'h31;
                    16'h994B: data_out = 8'h32;
                    16'h994C: data_out = 8'h33;
                    16'h994D: data_out = 8'h34;
                    16'h994E: data_out = 8'h35;
                    16'h994F: data_out = 8'h36;
                    16'h9950: data_out = 8'h37;
                    16'h9951: data_out = 8'h38;
                    16'h9952: data_out = 8'h39;
                    16'h9953: data_out = 8'h3A;
                    16'h9954: data_out = 8'h3B;
                    16'h9955: data_out = 8'h3C;
                    16'h9956: data_out = 8'h3D;
                    16'h9957: data_out = 8'h3E;
                    16'h9958: data_out = 8'h3F;
                    16'h9959: data_out = 8'h40;
                    16'h995A: data_out = 8'h41;
                    16'h995B: data_out = 8'h42;
                    16'h995C: data_out = 8'h43;
                    16'h995D: data_out = 8'h44;
                    16'h995E: data_out = 8'h45;
                    16'h995F: data_out = 8'h46;
                    16'h9960: data_out = 8'h47;
                    16'h9961: data_out = 8'h48;
                    16'h9962: data_out = 8'h49;
                    16'h9963: data_out = 8'h4A;
                    16'h9964: data_out = 8'h4B;
                    16'h9965: data_out = 8'h4C;
                    16'h9966: data_out = 8'h4D;
                    16'h9967: data_out = 8'h4E;
                    16'h9968: data_out = 8'h4F;
                    16'h9969: data_out = 8'h50;
                    16'h996A: data_out = 8'h51;
                    16'h996B: data_out = 8'h52;
                    16'h996C: data_out = 8'h53;
                    16'h996D: data_out = 8'h54;
                    16'h996E: data_out = 8'h55;
                    16'h996F: data_out = 8'h56;
                    16'h9970: data_out = 8'h57;
                    16'h9971: data_out = 8'h58;
                    16'h9972: data_out = 8'h59;
                    16'h9973: data_out = 8'h5A;
                    16'h9974: data_out = 8'h5B;
                    16'h9975: data_out = 8'h5C;
                    16'h9976: data_out = 8'h5D;
                    16'h9977: data_out = 8'h5E;
                    16'h9978: data_out = 8'h5F;
                    16'h9979: data_out = 8'h60;
                    16'h997A: data_out = 8'h61;
                    16'h997B: data_out = 8'h62;
                    16'h997C: data_out = 8'h63;
                    16'h997D: data_out = 8'h64;
                    16'h997E: data_out = 8'h65;
                    16'h997F: data_out = 8'h66;
                    16'h9980: data_out = 8'h99;
                    16'h9981: data_out = 8'h9A;
                    16'h9982: data_out = 8'h9B;
                    16'h9983: data_out = 8'h9C;
                    16'h9984: data_out = 8'h9D;
                    16'h9985: data_out = 8'h9E;
                    16'h9986: data_out = 8'h9F;
                    16'h9987: data_out = 8'hA0;
                    16'h9988: data_out = 8'hA1;
                    16'h9989: data_out = 8'hA2;
                    16'h998A: data_out = 8'hA3;
                    16'h998B: data_out = 8'hA4;
                    16'h998C: data_out = 8'hA5;
                    16'h998D: data_out = 8'hA6;
                    16'h998E: data_out = 8'hA7;
                    16'h998F: data_out = 8'hA8;
                    16'h9990: data_out = 8'hA9;
                    16'h9991: data_out = 8'hAA;
                    16'h9992: data_out = 8'hAB;
                    16'h9993: data_out = 8'hAC;
                    16'h9994: data_out = 8'hAD;
                    16'h9995: data_out = 8'hAE;
                    16'h9996: data_out = 8'hAF;
                    16'h9997: data_out = 8'hB0;
                    16'h9998: data_out = 8'hB1;
                    16'h9999: data_out = 8'hB2;
                    16'h999A: data_out = 8'hB3;
                    16'h999B: data_out = 8'hB4;
                    16'h999C: data_out = 8'hB5;
                    16'h999D: data_out = 8'hB6;
                    16'h999E: data_out = 8'hB7;
                    16'h999F: data_out = 8'hB8;
                    16'h99A0: data_out = 8'hB9;
                    16'h99A1: data_out = 8'hBA;
                    16'h99A2: data_out = 8'hBB;
                    16'h99A3: data_out = 8'hBC;
                    16'h99A4: data_out = 8'hBD;
                    16'h99A5: data_out = 8'hBE;
                    16'h99A6: data_out = 8'hBF;
                    16'h99A7: data_out = 8'hC0;
                    16'h99A8: data_out = 8'hC1;
                    16'h99A9: data_out = 8'hC2;
                    16'h99AA: data_out = 8'hC3;
                    16'h99AB: data_out = 8'hC4;
                    16'h99AC: data_out = 8'hC5;
                    16'h99AD: data_out = 8'hC6;
                    16'h99AE: data_out = 8'hC7;
                    16'h99AF: data_out = 8'hC8;
                    16'h99B0: data_out = 8'hC9;
                    16'h99B1: data_out = 8'hCA;
                    16'h99B2: data_out = 8'hCB;
                    16'h99B3: data_out = 8'hCC;
                    16'h99B4: data_out = 8'hCD;
                    16'h99B5: data_out = 8'hCE;
                    16'h99B6: data_out = 8'hCF;
                    16'h99B7: data_out = 8'hD0;
                    16'h99B8: data_out = 8'hD1;
                    16'h99B9: data_out = 8'hD2;
                    16'h99BA: data_out = 8'hD3;
                    16'h99BB: data_out = 8'hD4;
                    16'h99BC: data_out = 8'hD5;
                    16'h99BD: data_out = 8'hD6;
                    16'h99BE: data_out = 8'hD7;
                    16'h99BF: data_out = 8'hD8;
                    16'h99C0: data_out = 8'hD9;
                    16'h99C1: data_out = 8'hDA;
                    16'h99C2: data_out = 8'hDB;
                    16'h99C3: data_out = 8'hDC;
                    16'h99C4: data_out = 8'hDD;
                    16'h99C5: data_out = 8'hDE;
                    16'h99C6: data_out = 8'hDF;
                    16'h99C7: data_out = 8'hE0;
                    16'h99C8: data_out = 8'hE1;
                    16'h99C9: data_out = 8'hE2;
                    16'h99CA: data_out = 8'hE3;
                    16'h99CB: data_out = 8'hE4;
                    16'h99CC: data_out = 8'hE5;
                    16'h99CD: data_out = 8'hE6;
                    16'h99CE: data_out = 8'hE7;
                    16'h99CF: data_out = 8'hE8;
                    16'h99D0: data_out = 8'hE9;
                    16'h99D1: data_out = 8'hEA;
                    16'h99D2: data_out = 8'hEB;
                    16'h99D3: data_out = 8'hEC;
                    16'h99D4: data_out = 8'hED;
                    16'h99D5: data_out = 8'hEE;
                    16'h99D6: data_out = 8'hEF;
                    16'h99D7: data_out = 8'hF0;
                    16'h99D8: data_out = 8'hF1;
                    16'h99D9: data_out = 8'hF2;
                    16'h99DA: data_out = 8'hF3;
                    16'h99DB: data_out = 8'hF4;
                    16'h99DC: data_out = 8'hF5;
                    16'h99DD: data_out = 8'hF6;
                    16'h99DE: data_out = 8'hF7;
                    16'h99DF: data_out = 8'hF8;
                    16'h99E0: data_out = 8'hF9;
                    16'h99E1: data_out = 8'hFA;
                    16'h99E2: data_out = 8'hFB;
                    16'h99E3: data_out = 8'hFC;
                    16'h99E4: data_out = 8'hFD;
                    16'h99E5: data_out = 8'hFE;
                    16'h99E6: data_out = 8'hFF;
                    16'h99E7: data_out = 8'h80;
                    16'h99E8: data_out = 8'h81;
                    16'h99E9: data_out = 8'h82;
                    16'h99EA: data_out = 8'h83;
                    16'h99EB: data_out = 8'h84;
                    16'h99EC: data_out = 8'h85;
                    16'h99ED: data_out = 8'h86;
                    16'h99EE: data_out = 8'h87;
                    16'h99EF: data_out = 8'h88;
                    16'h99F0: data_out = 8'h89;
                    16'h99F1: data_out = 8'h8A;
                    16'h99F2: data_out = 8'h8B;
                    16'h99F3: data_out = 8'h8C;
                    16'h99F4: data_out = 8'h8D;
                    16'h99F5: data_out = 8'h8E;
                    16'h99F6: data_out = 8'h8F;
                    16'h99F7: data_out = 8'h90;
                    16'h99F8: data_out = 8'h91;
                    16'h99F9: data_out = 8'h92;
                    16'h99FA: data_out = 8'h93;
                    16'h99FB: data_out = 8'h94;
                    16'h99FC: data_out = 8'h95;
                    16'h99FD: data_out = 8'h96;
                    16'h99FE: data_out = 8'h97;
                    16'h99FF: data_out = 8'h98;
                    16'h9A00: data_out = 8'h9A;
                    16'h9A01: data_out = 8'h99;
                    16'h9A02: data_out = 8'h98;
                    16'h9A03: data_out = 8'h97;
                    16'h9A04: data_out = 8'h96;
                    16'h9A05: data_out = 8'h95;
                    16'h9A06: data_out = 8'h94;
                    16'h9A07: data_out = 8'h93;
                    16'h9A08: data_out = 8'h92;
                    16'h9A09: data_out = 8'h91;
                    16'h9A0A: data_out = 8'h90;
                    16'h9A0B: data_out = 8'h8F;
                    16'h9A0C: data_out = 8'h8E;
                    16'h9A0D: data_out = 8'h8D;
                    16'h9A0E: data_out = 8'h8C;
                    16'h9A0F: data_out = 8'h8B;
                    16'h9A10: data_out = 8'h8A;
                    16'h9A11: data_out = 8'h89;
                    16'h9A12: data_out = 8'h88;
                    16'h9A13: data_out = 8'h87;
                    16'h9A14: data_out = 8'h86;
                    16'h9A15: data_out = 8'h85;
                    16'h9A16: data_out = 8'h84;
                    16'h9A17: data_out = 8'h83;
                    16'h9A18: data_out = 8'h82;
                    16'h9A19: data_out = 8'h81;
                    16'h9A1A: data_out = 8'h0;
                    16'h9A1B: data_out = 8'h1;
                    16'h9A1C: data_out = 8'h2;
                    16'h9A1D: data_out = 8'h3;
                    16'h9A1E: data_out = 8'h4;
                    16'h9A1F: data_out = 8'h5;
                    16'h9A20: data_out = 8'h6;
                    16'h9A21: data_out = 8'h7;
                    16'h9A22: data_out = 8'h8;
                    16'h9A23: data_out = 8'h9;
                    16'h9A24: data_out = 8'hA;
                    16'h9A25: data_out = 8'hB;
                    16'h9A26: data_out = 8'hC;
                    16'h9A27: data_out = 8'hD;
                    16'h9A28: data_out = 8'hE;
                    16'h9A29: data_out = 8'hF;
                    16'h9A2A: data_out = 8'h10;
                    16'h9A2B: data_out = 8'h11;
                    16'h9A2C: data_out = 8'h12;
                    16'h9A2D: data_out = 8'h13;
                    16'h9A2E: data_out = 8'h14;
                    16'h9A2F: data_out = 8'h15;
                    16'h9A30: data_out = 8'h16;
                    16'h9A31: data_out = 8'h17;
                    16'h9A32: data_out = 8'h18;
                    16'h9A33: data_out = 8'h19;
                    16'h9A34: data_out = 8'h1A;
                    16'h9A35: data_out = 8'h1B;
                    16'h9A36: data_out = 8'h1C;
                    16'h9A37: data_out = 8'h1D;
                    16'h9A38: data_out = 8'h1E;
                    16'h9A39: data_out = 8'h1F;
                    16'h9A3A: data_out = 8'h20;
                    16'h9A3B: data_out = 8'h21;
                    16'h9A3C: data_out = 8'h22;
                    16'h9A3D: data_out = 8'h23;
                    16'h9A3E: data_out = 8'h24;
                    16'h9A3F: data_out = 8'h25;
                    16'h9A40: data_out = 8'h26;
                    16'h9A41: data_out = 8'h27;
                    16'h9A42: data_out = 8'h28;
                    16'h9A43: data_out = 8'h29;
                    16'h9A44: data_out = 8'h2A;
                    16'h9A45: data_out = 8'h2B;
                    16'h9A46: data_out = 8'h2C;
                    16'h9A47: data_out = 8'h2D;
                    16'h9A48: data_out = 8'h2E;
                    16'h9A49: data_out = 8'h2F;
                    16'h9A4A: data_out = 8'h30;
                    16'h9A4B: data_out = 8'h31;
                    16'h9A4C: data_out = 8'h32;
                    16'h9A4D: data_out = 8'h33;
                    16'h9A4E: data_out = 8'h34;
                    16'h9A4F: data_out = 8'h35;
                    16'h9A50: data_out = 8'h36;
                    16'h9A51: data_out = 8'h37;
                    16'h9A52: data_out = 8'h38;
                    16'h9A53: data_out = 8'h39;
                    16'h9A54: data_out = 8'h3A;
                    16'h9A55: data_out = 8'h3B;
                    16'h9A56: data_out = 8'h3C;
                    16'h9A57: data_out = 8'h3D;
                    16'h9A58: data_out = 8'h3E;
                    16'h9A59: data_out = 8'h3F;
                    16'h9A5A: data_out = 8'h40;
                    16'h9A5B: data_out = 8'h41;
                    16'h9A5C: data_out = 8'h42;
                    16'h9A5D: data_out = 8'h43;
                    16'h9A5E: data_out = 8'h44;
                    16'h9A5F: data_out = 8'h45;
                    16'h9A60: data_out = 8'h46;
                    16'h9A61: data_out = 8'h47;
                    16'h9A62: data_out = 8'h48;
                    16'h9A63: data_out = 8'h49;
                    16'h9A64: data_out = 8'h4A;
                    16'h9A65: data_out = 8'h4B;
                    16'h9A66: data_out = 8'h4C;
                    16'h9A67: data_out = 8'h4D;
                    16'h9A68: data_out = 8'h4E;
                    16'h9A69: data_out = 8'h4F;
                    16'h9A6A: data_out = 8'h50;
                    16'h9A6B: data_out = 8'h51;
                    16'h9A6C: data_out = 8'h52;
                    16'h9A6D: data_out = 8'h53;
                    16'h9A6E: data_out = 8'h54;
                    16'h9A6F: data_out = 8'h55;
                    16'h9A70: data_out = 8'h56;
                    16'h9A71: data_out = 8'h57;
                    16'h9A72: data_out = 8'h58;
                    16'h9A73: data_out = 8'h59;
                    16'h9A74: data_out = 8'h5A;
                    16'h9A75: data_out = 8'h5B;
                    16'h9A76: data_out = 8'h5C;
                    16'h9A77: data_out = 8'h5D;
                    16'h9A78: data_out = 8'h5E;
                    16'h9A79: data_out = 8'h5F;
                    16'h9A7A: data_out = 8'h60;
                    16'h9A7B: data_out = 8'h61;
                    16'h9A7C: data_out = 8'h62;
                    16'h9A7D: data_out = 8'h63;
                    16'h9A7E: data_out = 8'h64;
                    16'h9A7F: data_out = 8'h65;
                    16'h9A80: data_out = 8'h9A;
                    16'h9A81: data_out = 8'h9B;
                    16'h9A82: data_out = 8'h9C;
                    16'h9A83: data_out = 8'h9D;
                    16'h9A84: data_out = 8'h9E;
                    16'h9A85: data_out = 8'h9F;
                    16'h9A86: data_out = 8'hA0;
                    16'h9A87: data_out = 8'hA1;
                    16'h9A88: data_out = 8'hA2;
                    16'h9A89: data_out = 8'hA3;
                    16'h9A8A: data_out = 8'hA4;
                    16'h9A8B: data_out = 8'hA5;
                    16'h9A8C: data_out = 8'hA6;
                    16'h9A8D: data_out = 8'hA7;
                    16'h9A8E: data_out = 8'hA8;
                    16'h9A8F: data_out = 8'hA9;
                    16'h9A90: data_out = 8'hAA;
                    16'h9A91: data_out = 8'hAB;
                    16'h9A92: data_out = 8'hAC;
                    16'h9A93: data_out = 8'hAD;
                    16'h9A94: data_out = 8'hAE;
                    16'h9A95: data_out = 8'hAF;
                    16'h9A96: data_out = 8'hB0;
                    16'h9A97: data_out = 8'hB1;
                    16'h9A98: data_out = 8'hB2;
                    16'h9A99: data_out = 8'hB3;
                    16'h9A9A: data_out = 8'hB4;
                    16'h9A9B: data_out = 8'hB5;
                    16'h9A9C: data_out = 8'hB6;
                    16'h9A9D: data_out = 8'hB7;
                    16'h9A9E: data_out = 8'hB8;
                    16'h9A9F: data_out = 8'hB9;
                    16'h9AA0: data_out = 8'hBA;
                    16'h9AA1: data_out = 8'hBB;
                    16'h9AA2: data_out = 8'hBC;
                    16'h9AA3: data_out = 8'hBD;
                    16'h9AA4: data_out = 8'hBE;
                    16'h9AA5: data_out = 8'hBF;
                    16'h9AA6: data_out = 8'hC0;
                    16'h9AA7: data_out = 8'hC1;
                    16'h9AA8: data_out = 8'hC2;
                    16'h9AA9: data_out = 8'hC3;
                    16'h9AAA: data_out = 8'hC4;
                    16'h9AAB: data_out = 8'hC5;
                    16'h9AAC: data_out = 8'hC6;
                    16'h9AAD: data_out = 8'hC7;
                    16'h9AAE: data_out = 8'hC8;
                    16'h9AAF: data_out = 8'hC9;
                    16'h9AB0: data_out = 8'hCA;
                    16'h9AB1: data_out = 8'hCB;
                    16'h9AB2: data_out = 8'hCC;
                    16'h9AB3: data_out = 8'hCD;
                    16'h9AB4: data_out = 8'hCE;
                    16'h9AB5: data_out = 8'hCF;
                    16'h9AB6: data_out = 8'hD0;
                    16'h9AB7: data_out = 8'hD1;
                    16'h9AB8: data_out = 8'hD2;
                    16'h9AB9: data_out = 8'hD3;
                    16'h9ABA: data_out = 8'hD4;
                    16'h9ABB: data_out = 8'hD5;
                    16'h9ABC: data_out = 8'hD6;
                    16'h9ABD: data_out = 8'hD7;
                    16'h9ABE: data_out = 8'hD8;
                    16'h9ABF: data_out = 8'hD9;
                    16'h9AC0: data_out = 8'hDA;
                    16'h9AC1: data_out = 8'hDB;
                    16'h9AC2: data_out = 8'hDC;
                    16'h9AC3: data_out = 8'hDD;
                    16'h9AC4: data_out = 8'hDE;
                    16'h9AC5: data_out = 8'hDF;
                    16'h9AC6: data_out = 8'hE0;
                    16'h9AC7: data_out = 8'hE1;
                    16'h9AC8: data_out = 8'hE2;
                    16'h9AC9: data_out = 8'hE3;
                    16'h9ACA: data_out = 8'hE4;
                    16'h9ACB: data_out = 8'hE5;
                    16'h9ACC: data_out = 8'hE6;
                    16'h9ACD: data_out = 8'hE7;
                    16'h9ACE: data_out = 8'hE8;
                    16'h9ACF: data_out = 8'hE9;
                    16'h9AD0: data_out = 8'hEA;
                    16'h9AD1: data_out = 8'hEB;
                    16'h9AD2: data_out = 8'hEC;
                    16'h9AD3: data_out = 8'hED;
                    16'h9AD4: data_out = 8'hEE;
                    16'h9AD5: data_out = 8'hEF;
                    16'h9AD6: data_out = 8'hF0;
                    16'h9AD7: data_out = 8'hF1;
                    16'h9AD8: data_out = 8'hF2;
                    16'h9AD9: data_out = 8'hF3;
                    16'h9ADA: data_out = 8'hF4;
                    16'h9ADB: data_out = 8'hF5;
                    16'h9ADC: data_out = 8'hF6;
                    16'h9ADD: data_out = 8'hF7;
                    16'h9ADE: data_out = 8'hF8;
                    16'h9ADF: data_out = 8'hF9;
                    16'h9AE0: data_out = 8'hFA;
                    16'h9AE1: data_out = 8'hFB;
                    16'h9AE2: data_out = 8'hFC;
                    16'h9AE3: data_out = 8'hFD;
                    16'h9AE4: data_out = 8'hFE;
                    16'h9AE5: data_out = 8'hFF;
                    16'h9AE6: data_out = 8'h80;
                    16'h9AE7: data_out = 8'h81;
                    16'h9AE8: data_out = 8'h82;
                    16'h9AE9: data_out = 8'h83;
                    16'h9AEA: data_out = 8'h84;
                    16'h9AEB: data_out = 8'h85;
                    16'h9AEC: data_out = 8'h86;
                    16'h9AED: data_out = 8'h87;
                    16'h9AEE: data_out = 8'h88;
                    16'h9AEF: data_out = 8'h89;
                    16'h9AF0: data_out = 8'h8A;
                    16'h9AF1: data_out = 8'h8B;
                    16'h9AF2: data_out = 8'h8C;
                    16'h9AF3: data_out = 8'h8D;
                    16'h9AF4: data_out = 8'h8E;
                    16'h9AF5: data_out = 8'h8F;
                    16'h9AF6: data_out = 8'h90;
                    16'h9AF7: data_out = 8'h91;
                    16'h9AF8: data_out = 8'h92;
                    16'h9AF9: data_out = 8'h93;
                    16'h9AFA: data_out = 8'h94;
                    16'h9AFB: data_out = 8'h95;
                    16'h9AFC: data_out = 8'h96;
                    16'h9AFD: data_out = 8'h97;
                    16'h9AFE: data_out = 8'h98;
                    16'h9AFF: data_out = 8'h99;
                    16'h9B00: data_out = 8'h9B;
                    16'h9B01: data_out = 8'h9A;
                    16'h9B02: data_out = 8'h99;
                    16'h9B03: data_out = 8'h98;
                    16'h9B04: data_out = 8'h97;
                    16'h9B05: data_out = 8'h96;
                    16'h9B06: data_out = 8'h95;
                    16'h9B07: data_out = 8'h94;
                    16'h9B08: data_out = 8'h93;
                    16'h9B09: data_out = 8'h92;
                    16'h9B0A: data_out = 8'h91;
                    16'h9B0B: data_out = 8'h90;
                    16'h9B0C: data_out = 8'h8F;
                    16'h9B0D: data_out = 8'h8E;
                    16'h9B0E: data_out = 8'h8D;
                    16'h9B0F: data_out = 8'h8C;
                    16'h9B10: data_out = 8'h8B;
                    16'h9B11: data_out = 8'h8A;
                    16'h9B12: data_out = 8'h89;
                    16'h9B13: data_out = 8'h88;
                    16'h9B14: data_out = 8'h87;
                    16'h9B15: data_out = 8'h86;
                    16'h9B16: data_out = 8'h85;
                    16'h9B17: data_out = 8'h84;
                    16'h9B18: data_out = 8'h83;
                    16'h9B19: data_out = 8'h82;
                    16'h9B1A: data_out = 8'h81;
                    16'h9B1B: data_out = 8'h0;
                    16'h9B1C: data_out = 8'h1;
                    16'h9B1D: data_out = 8'h2;
                    16'h9B1E: data_out = 8'h3;
                    16'h9B1F: data_out = 8'h4;
                    16'h9B20: data_out = 8'h5;
                    16'h9B21: data_out = 8'h6;
                    16'h9B22: data_out = 8'h7;
                    16'h9B23: data_out = 8'h8;
                    16'h9B24: data_out = 8'h9;
                    16'h9B25: data_out = 8'hA;
                    16'h9B26: data_out = 8'hB;
                    16'h9B27: data_out = 8'hC;
                    16'h9B28: data_out = 8'hD;
                    16'h9B29: data_out = 8'hE;
                    16'h9B2A: data_out = 8'hF;
                    16'h9B2B: data_out = 8'h10;
                    16'h9B2C: data_out = 8'h11;
                    16'h9B2D: data_out = 8'h12;
                    16'h9B2E: data_out = 8'h13;
                    16'h9B2F: data_out = 8'h14;
                    16'h9B30: data_out = 8'h15;
                    16'h9B31: data_out = 8'h16;
                    16'h9B32: data_out = 8'h17;
                    16'h9B33: data_out = 8'h18;
                    16'h9B34: data_out = 8'h19;
                    16'h9B35: data_out = 8'h1A;
                    16'h9B36: data_out = 8'h1B;
                    16'h9B37: data_out = 8'h1C;
                    16'h9B38: data_out = 8'h1D;
                    16'h9B39: data_out = 8'h1E;
                    16'h9B3A: data_out = 8'h1F;
                    16'h9B3B: data_out = 8'h20;
                    16'h9B3C: data_out = 8'h21;
                    16'h9B3D: data_out = 8'h22;
                    16'h9B3E: data_out = 8'h23;
                    16'h9B3F: data_out = 8'h24;
                    16'h9B40: data_out = 8'h25;
                    16'h9B41: data_out = 8'h26;
                    16'h9B42: data_out = 8'h27;
                    16'h9B43: data_out = 8'h28;
                    16'h9B44: data_out = 8'h29;
                    16'h9B45: data_out = 8'h2A;
                    16'h9B46: data_out = 8'h2B;
                    16'h9B47: data_out = 8'h2C;
                    16'h9B48: data_out = 8'h2D;
                    16'h9B49: data_out = 8'h2E;
                    16'h9B4A: data_out = 8'h2F;
                    16'h9B4B: data_out = 8'h30;
                    16'h9B4C: data_out = 8'h31;
                    16'h9B4D: data_out = 8'h32;
                    16'h9B4E: data_out = 8'h33;
                    16'h9B4F: data_out = 8'h34;
                    16'h9B50: data_out = 8'h35;
                    16'h9B51: data_out = 8'h36;
                    16'h9B52: data_out = 8'h37;
                    16'h9B53: data_out = 8'h38;
                    16'h9B54: data_out = 8'h39;
                    16'h9B55: data_out = 8'h3A;
                    16'h9B56: data_out = 8'h3B;
                    16'h9B57: data_out = 8'h3C;
                    16'h9B58: data_out = 8'h3D;
                    16'h9B59: data_out = 8'h3E;
                    16'h9B5A: data_out = 8'h3F;
                    16'h9B5B: data_out = 8'h40;
                    16'h9B5C: data_out = 8'h41;
                    16'h9B5D: data_out = 8'h42;
                    16'h9B5E: data_out = 8'h43;
                    16'h9B5F: data_out = 8'h44;
                    16'h9B60: data_out = 8'h45;
                    16'h9B61: data_out = 8'h46;
                    16'h9B62: data_out = 8'h47;
                    16'h9B63: data_out = 8'h48;
                    16'h9B64: data_out = 8'h49;
                    16'h9B65: data_out = 8'h4A;
                    16'h9B66: data_out = 8'h4B;
                    16'h9B67: data_out = 8'h4C;
                    16'h9B68: data_out = 8'h4D;
                    16'h9B69: data_out = 8'h4E;
                    16'h9B6A: data_out = 8'h4F;
                    16'h9B6B: data_out = 8'h50;
                    16'h9B6C: data_out = 8'h51;
                    16'h9B6D: data_out = 8'h52;
                    16'h9B6E: data_out = 8'h53;
                    16'h9B6F: data_out = 8'h54;
                    16'h9B70: data_out = 8'h55;
                    16'h9B71: data_out = 8'h56;
                    16'h9B72: data_out = 8'h57;
                    16'h9B73: data_out = 8'h58;
                    16'h9B74: data_out = 8'h59;
                    16'h9B75: data_out = 8'h5A;
                    16'h9B76: data_out = 8'h5B;
                    16'h9B77: data_out = 8'h5C;
                    16'h9B78: data_out = 8'h5D;
                    16'h9B79: data_out = 8'h5E;
                    16'h9B7A: data_out = 8'h5F;
                    16'h9B7B: data_out = 8'h60;
                    16'h9B7C: data_out = 8'h61;
                    16'h9B7D: data_out = 8'h62;
                    16'h9B7E: data_out = 8'h63;
                    16'h9B7F: data_out = 8'h64;
                    16'h9B80: data_out = 8'h9B;
                    16'h9B81: data_out = 8'h9C;
                    16'h9B82: data_out = 8'h9D;
                    16'h9B83: data_out = 8'h9E;
                    16'h9B84: data_out = 8'h9F;
                    16'h9B85: data_out = 8'hA0;
                    16'h9B86: data_out = 8'hA1;
                    16'h9B87: data_out = 8'hA2;
                    16'h9B88: data_out = 8'hA3;
                    16'h9B89: data_out = 8'hA4;
                    16'h9B8A: data_out = 8'hA5;
                    16'h9B8B: data_out = 8'hA6;
                    16'h9B8C: data_out = 8'hA7;
                    16'h9B8D: data_out = 8'hA8;
                    16'h9B8E: data_out = 8'hA9;
                    16'h9B8F: data_out = 8'hAA;
                    16'h9B90: data_out = 8'hAB;
                    16'h9B91: data_out = 8'hAC;
                    16'h9B92: data_out = 8'hAD;
                    16'h9B93: data_out = 8'hAE;
                    16'h9B94: data_out = 8'hAF;
                    16'h9B95: data_out = 8'hB0;
                    16'h9B96: data_out = 8'hB1;
                    16'h9B97: data_out = 8'hB2;
                    16'h9B98: data_out = 8'hB3;
                    16'h9B99: data_out = 8'hB4;
                    16'h9B9A: data_out = 8'hB5;
                    16'h9B9B: data_out = 8'hB6;
                    16'h9B9C: data_out = 8'hB7;
                    16'h9B9D: data_out = 8'hB8;
                    16'h9B9E: data_out = 8'hB9;
                    16'h9B9F: data_out = 8'hBA;
                    16'h9BA0: data_out = 8'hBB;
                    16'h9BA1: data_out = 8'hBC;
                    16'h9BA2: data_out = 8'hBD;
                    16'h9BA3: data_out = 8'hBE;
                    16'h9BA4: data_out = 8'hBF;
                    16'h9BA5: data_out = 8'hC0;
                    16'h9BA6: data_out = 8'hC1;
                    16'h9BA7: data_out = 8'hC2;
                    16'h9BA8: data_out = 8'hC3;
                    16'h9BA9: data_out = 8'hC4;
                    16'h9BAA: data_out = 8'hC5;
                    16'h9BAB: data_out = 8'hC6;
                    16'h9BAC: data_out = 8'hC7;
                    16'h9BAD: data_out = 8'hC8;
                    16'h9BAE: data_out = 8'hC9;
                    16'h9BAF: data_out = 8'hCA;
                    16'h9BB0: data_out = 8'hCB;
                    16'h9BB1: data_out = 8'hCC;
                    16'h9BB2: data_out = 8'hCD;
                    16'h9BB3: data_out = 8'hCE;
                    16'h9BB4: data_out = 8'hCF;
                    16'h9BB5: data_out = 8'hD0;
                    16'h9BB6: data_out = 8'hD1;
                    16'h9BB7: data_out = 8'hD2;
                    16'h9BB8: data_out = 8'hD3;
                    16'h9BB9: data_out = 8'hD4;
                    16'h9BBA: data_out = 8'hD5;
                    16'h9BBB: data_out = 8'hD6;
                    16'h9BBC: data_out = 8'hD7;
                    16'h9BBD: data_out = 8'hD8;
                    16'h9BBE: data_out = 8'hD9;
                    16'h9BBF: data_out = 8'hDA;
                    16'h9BC0: data_out = 8'hDB;
                    16'h9BC1: data_out = 8'hDC;
                    16'h9BC2: data_out = 8'hDD;
                    16'h9BC3: data_out = 8'hDE;
                    16'h9BC4: data_out = 8'hDF;
                    16'h9BC5: data_out = 8'hE0;
                    16'h9BC6: data_out = 8'hE1;
                    16'h9BC7: data_out = 8'hE2;
                    16'h9BC8: data_out = 8'hE3;
                    16'h9BC9: data_out = 8'hE4;
                    16'h9BCA: data_out = 8'hE5;
                    16'h9BCB: data_out = 8'hE6;
                    16'h9BCC: data_out = 8'hE7;
                    16'h9BCD: data_out = 8'hE8;
                    16'h9BCE: data_out = 8'hE9;
                    16'h9BCF: data_out = 8'hEA;
                    16'h9BD0: data_out = 8'hEB;
                    16'h9BD1: data_out = 8'hEC;
                    16'h9BD2: data_out = 8'hED;
                    16'h9BD3: data_out = 8'hEE;
                    16'h9BD4: data_out = 8'hEF;
                    16'h9BD5: data_out = 8'hF0;
                    16'h9BD6: data_out = 8'hF1;
                    16'h9BD7: data_out = 8'hF2;
                    16'h9BD8: data_out = 8'hF3;
                    16'h9BD9: data_out = 8'hF4;
                    16'h9BDA: data_out = 8'hF5;
                    16'h9BDB: data_out = 8'hF6;
                    16'h9BDC: data_out = 8'hF7;
                    16'h9BDD: data_out = 8'hF8;
                    16'h9BDE: data_out = 8'hF9;
                    16'h9BDF: data_out = 8'hFA;
                    16'h9BE0: data_out = 8'hFB;
                    16'h9BE1: data_out = 8'hFC;
                    16'h9BE2: data_out = 8'hFD;
                    16'h9BE3: data_out = 8'hFE;
                    16'h9BE4: data_out = 8'hFF;
                    16'h9BE5: data_out = 8'h80;
                    16'h9BE6: data_out = 8'h81;
                    16'h9BE7: data_out = 8'h82;
                    16'h9BE8: data_out = 8'h83;
                    16'h9BE9: data_out = 8'h84;
                    16'h9BEA: data_out = 8'h85;
                    16'h9BEB: data_out = 8'h86;
                    16'h9BEC: data_out = 8'h87;
                    16'h9BED: data_out = 8'h88;
                    16'h9BEE: data_out = 8'h89;
                    16'h9BEF: data_out = 8'h8A;
                    16'h9BF0: data_out = 8'h8B;
                    16'h9BF1: data_out = 8'h8C;
                    16'h9BF2: data_out = 8'h8D;
                    16'h9BF3: data_out = 8'h8E;
                    16'h9BF4: data_out = 8'h8F;
                    16'h9BF5: data_out = 8'h90;
                    16'h9BF6: data_out = 8'h91;
                    16'h9BF7: data_out = 8'h92;
                    16'h9BF8: data_out = 8'h93;
                    16'h9BF9: data_out = 8'h94;
                    16'h9BFA: data_out = 8'h95;
                    16'h9BFB: data_out = 8'h96;
                    16'h9BFC: data_out = 8'h97;
                    16'h9BFD: data_out = 8'h98;
                    16'h9BFE: data_out = 8'h99;
                    16'h9BFF: data_out = 8'h9A;
                    16'h9C00: data_out = 8'h9C;
                    16'h9C01: data_out = 8'h9B;
                    16'h9C02: data_out = 8'h9A;
                    16'h9C03: data_out = 8'h99;
                    16'h9C04: data_out = 8'h98;
                    16'h9C05: data_out = 8'h97;
                    16'h9C06: data_out = 8'h96;
                    16'h9C07: data_out = 8'h95;
                    16'h9C08: data_out = 8'h94;
                    16'h9C09: data_out = 8'h93;
                    16'h9C0A: data_out = 8'h92;
                    16'h9C0B: data_out = 8'h91;
                    16'h9C0C: data_out = 8'h90;
                    16'h9C0D: data_out = 8'h8F;
                    16'h9C0E: data_out = 8'h8E;
                    16'h9C0F: data_out = 8'h8D;
                    16'h9C10: data_out = 8'h8C;
                    16'h9C11: data_out = 8'h8B;
                    16'h9C12: data_out = 8'h8A;
                    16'h9C13: data_out = 8'h89;
                    16'h9C14: data_out = 8'h88;
                    16'h9C15: data_out = 8'h87;
                    16'h9C16: data_out = 8'h86;
                    16'h9C17: data_out = 8'h85;
                    16'h9C18: data_out = 8'h84;
                    16'h9C19: data_out = 8'h83;
                    16'h9C1A: data_out = 8'h82;
                    16'h9C1B: data_out = 8'h81;
                    16'h9C1C: data_out = 8'h0;
                    16'h9C1D: data_out = 8'h1;
                    16'h9C1E: data_out = 8'h2;
                    16'h9C1F: data_out = 8'h3;
                    16'h9C20: data_out = 8'h4;
                    16'h9C21: data_out = 8'h5;
                    16'h9C22: data_out = 8'h6;
                    16'h9C23: data_out = 8'h7;
                    16'h9C24: data_out = 8'h8;
                    16'h9C25: data_out = 8'h9;
                    16'h9C26: data_out = 8'hA;
                    16'h9C27: data_out = 8'hB;
                    16'h9C28: data_out = 8'hC;
                    16'h9C29: data_out = 8'hD;
                    16'h9C2A: data_out = 8'hE;
                    16'h9C2B: data_out = 8'hF;
                    16'h9C2C: data_out = 8'h10;
                    16'h9C2D: data_out = 8'h11;
                    16'h9C2E: data_out = 8'h12;
                    16'h9C2F: data_out = 8'h13;
                    16'h9C30: data_out = 8'h14;
                    16'h9C31: data_out = 8'h15;
                    16'h9C32: data_out = 8'h16;
                    16'h9C33: data_out = 8'h17;
                    16'h9C34: data_out = 8'h18;
                    16'h9C35: data_out = 8'h19;
                    16'h9C36: data_out = 8'h1A;
                    16'h9C37: data_out = 8'h1B;
                    16'h9C38: data_out = 8'h1C;
                    16'h9C39: data_out = 8'h1D;
                    16'h9C3A: data_out = 8'h1E;
                    16'h9C3B: data_out = 8'h1F;
                    16'h9C3C: data_out = 8'h20;
                    16'h9C3D: data_out = 8'h21;
                    16'h9C3E: data_out = 8'h22;
                    16'h9C3F: data_out = 8'h23;
                    16'h9C40: data_out = 8'h24;
                    16'h9C41: data_out = 8'h25;
                    16'h9C42: data_out = 8'h26;
                    16'h9C43: data_out = 8'h27;
                    16'h9C44: data_out = 8'h28;
                    16'h9C45: data_out = 8'h29;
                    16'h9C46: data_out = 8'h2A;
                    16'h9C47: data_out = 8'h2B;
                    16'h9C48: data_out = 8'h2C;
                    16'h9C49: data_out = 8'h2D;
                    16'h9C4A: data_out = 8'h2E;
                    16'h9C4B: data_out = 8'h2F;
                    16'h9C4C: data_out = 8'h30;
                    16'h9C4D: data_out = 8'h31;
                    16'h9C4E: data_out = 8'h32;
                    16'h9C4F: data_out = 8'h33;
                    16'h9C50: data_out = 8'h34;
                    16'h9C51: data_out = 8'h35;
                    16'h9C52: data_out = 8'h36;
                    16'h9C53: data_out = 8'h37;
                    16'h9C54: data_out = 8'h38;
                    16'h9C55: data_out = 8'h39;
                    16'h9C56: data_out = 8'h3A;
                    16'h9C57: data_out = 8'h3B;
                    16'h9C58: data_out = 8'h3C;
                    16'h9C59: data_out = 8'h3D;
                    16'h9C5A: data_out = 8'h3E;
                    16'h9C5B: data_out = 8'h3F;
                    16'h9C5C: data_out = 8'h40;
                    16'h9C5D: data_out = 8'h41;
                    16'h9C5E: data_out = 8'h42;
                    16'h9C5F: data_out = 8'h43;
                    16'h9C60: data_out = 8'h44;
                    16'h9C61: data_out = 8'h45;
                    16'h9C62: data_out = 8'h46;
                    16'h9C63: data_out = 8'h47;
                    16'h9C64: data_out = 8'h48;
                    16'h9C65: data_out = 8'h49;
                    16'h9C66: data_out = 8'h4A;
                    16'h9C67: data_out = 8'h4B;
                    16'h9C68: data_out = 8'h4C;
                    16'h9C69: data_out = 8'h4D;
                    16'h9C6A: data_out = 8'h4E;
                    16'h9C6B: data_out = 8'h4F;
                    16'h9C6C: data_out = 8'h50;
                    16'h9C6D: data_out = 8'h51;
                    16'h9C6E: data_out = 8'h52;
                    16'h9C6F: data_out = 8'h53;
                    16'h9C70: data_out = 8'h54;
                    16'h9C71: data_out = 8'h55;
                    16'h9C72: data_out = 8'h56;
                    16'h9C73: data_out = 8'h57;
                    16'h9C74: data_out = 8'h58;
                    16'h9C75: data_out = 8'h59;
                    16'h9C76: data_out = 8'h5A;
                    16'h9C77: data_out = 8'h5B;
                    16'h9C78: data_out = 8'h5C;
                    16'h9C79: data_out = 8'h5D;
                    16'h9C7A: data_out = 8'h5E;
                    16'h9C7B: data_out = 8'h5F;
                    16'h9C7C: data_out = 8'h60;
                    16'h9C7D: data_out = 8'h61;
                    16'h9C7E: data_out = 8'h62;
                    16'h9C7F: data_out = 8'h63;
                    16'h9C80: data_out = 8'h9C;
                    16'h9C81: data_out = 8'h9D;
                    16'h9C82: data_out = 8'h9E;
                    16'h9C83: data_out = 8'h9F;
                    16'h9C84: data_out = 8'hA0;
                    16'h9C85: data_out = 8'hA1;
                    16'h9C86: data_out = 8'hA2;
                    16'h9C87: data_out = 8'hA3;
                    16'h9C88: data_out = 8'hA4;
                    16'h9C89: data_out = 8'hA5;
                    16'h9C8A: data_out = 8'hA6;
                    16'h9C8B: data_out = 8'hA7;
                    16'h9C8C: data_out = 8'hA8;
                    16'h9C8D: data_out = 8'hA9;
                    16'h9C8E: data_out = 8'hAA;
                    16'h9C8F: data_out = 8'hAB;
                    16'h9C90: data_out = 8'hAC;
                    16'h9C91: data_out = 8'hAD;
                    16'h9C92: data_out = 8'hAE;
                    16'h9C93: data_out = 8'hAF;
                    16'h9C94: data_out = 8'hB0;
                    16'h9C95: data_out = 8'hB1;
                    16'h9C96: data_out = 8'hB2;
                    16'h9C97: data_out = 8'hB3;
                    16'h9C98: data_out = 8'hB4;
                    16'h9C99: data_out = 8'hB5;
                    16'h9C9A: data_out = 8'hB6;
                    16'h9C9B: data_out = 8'hB7;
                    16'h9C9C: data_out = 8'hB8;
                    16'h9C9D: data_out = 8'hB9;
                    16'h9C9E: data_out = 8'hBA;
                    16'h9C9F: data_out = 8'hBB;
                    16'h9CA0: data_out = 8'hBC;
                    16'h9CA1: data_out = 8'hBD;
                    16'h9CA2: data_out = 8'hBE;
                    16'h9CA3: data_out = 8'hBF;
                    16'h9CA4: data_out = 8'hC0;
                    16'h9CA5: data_out = 8'hC1;
                    16'h9CA6: data_out = 8'hC2;
                    16'h9CA7: data_out = 8'hC3;
                    16'h9CA8: data_out = 8'hC4;
                    16'h9CA9: data_out = 8'hC5;
                    16'h9CAA: data_out = 8'hC6;
                    16'h9CAB: data_out = 8'hC7;
                    16'h9CAC: data_out = 8'hC8;
                    16'h9CAD: data_out = 8'hC9;
                    16'h9CAE: data_out = 8'hCA;
                    16'h9CAF: data_out = 8'hCB;
                    16'h9CB0: data_out = 8'hCC;
                    16'h9CB1: data_out = 8'hCD;
                    16'h9CB2: data_out = 8'hCE;
                    16'h9CB3: data_out = 8'hCF;
                    16'h9CB4: data_out = 8'hD0;
                    16'h9CB5: data_out = 8'hD1;
                    16'h9CB6: data_out = 8'hD2;
                    16'h9CB7: data_out = 8'hD3;
                    16'h9CB8: data_out = 8'hD4;
                    16'h9CB9: data_out = 8'hD5;
                    16'h9CBA: data_out = 8'hD6;
                    16'h9CBB: data_out = 8'hD7;
                    16'h9CBC: data_out = 8'hD8;
                    16'h9CBD: data_out = 8'hD9;
                    16'h9CBE: data_out = 8'hDA;
                    16'h9CBF: data_out = 8'hDB;
                    16'h9CC0: data_out = 8'hDC;
                    16'h9CC1: data_out = 8'hDD;
                    16'h9CC2: data_out = 8'hDE;
                    16'h9CC3: data_out = 8'hDF;
                    16'h9CC4: data_out = 8'hE0;
                    16'h9CC5: data_out = 8'hE1;
                    16'h9CC6: data_out = 8'hE2;
                    16'h9CC7: data_out = 8'hE3;
                    16'h9CC8: data_out = 8'hE4;
                    16'h9CC9: data_out = 8'hE5;
                    16'h9CCA: data_out = 8'hE6;
                    16'h9CCB: data_out = 8'hE7;
                    16'h9CCC: data_out = 8'hE8;
                    16'h9CCD: data_out = 8'hE9;
                    16'h9CCE: data_out = 8'hEA;
                    16'h9CCF: data_out = 8'hEB;
                    16'h9CD0: data_out = 8'hEC;
                    16'h9CD1: data_out = 8'hED;
                    16'h9CD2: data_out = 8'hEE;
                    16'h9CD3: data_out = 8'hEF;
                    16'h9CD4: data_out = 8'hF0;
                    16'h9CD5: data_out = 8'hF1;
                    16'h9CD6: data_out = 8'hF2;
                    16'h9CD7: data_out = 8'hF3;
                    16'h9CD8: data_out = 8'hF4;
                    16'h9CD9: data_out = 8'hF5;
                    16'h9CDA: data_out = 8'hF6;
                    16'h9CDB: data_out = 8'hF7;
                    16'h9CDC: data_out = 8'hF8;
                    16'h9CDD: data_out = 8'hF9;
                    16'h9CDE: data_out = 8'hFA;
                    16'h9CDF: data_out = 8'hFB;
                    16'h9CE0: data_out = 8'hFC;
                    16'h9CE1: data_out = 8'hFD;
                    16'h9CE2: data_out = 8'hFE;
                    16'h9CE3: data_out = 8'hFF;
                    16'h9CE4: data_out = 8'h80;
                    16'h9CE5: data_out = 8'h81;
                    16'h9CE6: data_out = 8'h82;
                    16'h9CE7: data_out = 8'h83;
                    16'h9CE8: data_out = 8'h84;
                    16'h9CE9: data_out = 8'h85;
                    16'h9CEA: data_out = 8'h86;
                    16'h9CEB: data_out = 8'h87;
                    16'h9CEC: data_out = 8'h88;
                    16'h9CED: data_out = 8'h89;
                    16'h9CEE: data_out = 8'h8A;
                    16'h9CEF: data_out = 8'h8B;
                    16'h9CF0: data_out = 8'h8C;
                    16'h9CF1: data_out = 8'h8D;
                    16'h9CF2: data_out = 8'h8E;
                    16'h9CF3: data_out = 8'h8F;
                    16'h9CF4: data_out = 8'h90;
                    16'h9CF5: data_out = 8'h91;
                    16'h9CF6: data_out = 8'h92;
                    16'h9CF7: data_out = 8'h93;
                    16'h9CF8: data_out = 8'h94;
                    16'h9CF9: data_out = 8'h95;
                    16'h9CFA: data_out = 8'h96;
                    16'h9CFB: data_out = 8'h97;
                    16'h9CFC: data_out = 8'h98;
                    16'h9CFD: data_out = 8'h99;
                    16'h9CFE: data_out = 8'h9A;
                    16'h9CFF: data_out = 8'h9B;
                    16'h9D00: data_out = 8'h9D;
                    16'h9D01: data_out = 8'h9C;
                    16'h9D02: data_out = 8'h9B;
                    16'h9D03: data_out = 8'h9A;
                    16'h9D04: data_out = 8'h99;
                    16'h9D05: data_out = 8'h98;
                    16'h9D06: data_out = 8'h97;
                    16'h9D07: data_out = 8'h96;
                    16'h9D08: data_out = 8'h95;
                    16'h9D09: data_out = 8'h94;
                    16'h9D0A: data_out = 8'h93;
                    16'h9D0B: data_out = 8'h92;
                    16'h9D0C: data_out = 8'h91;
                    16'h9D0D: data_out = 8'h90;
                    16'h9D0E: data_out = 8'h8F;
                    16'h9D0F: data_out = 8'h8E;
                    16'h9D10: data_out = 8'h8D;
                    16'h9D11: data_out = 8'h8C;
                    16'h9D12: data_out = 8'h8B;
                    16'h9D13: data_out = 8'h8A;
                    16'h9D14: data_out = 8'h89;
                    16'h9D15: data_out = 8'h88;
                    16'h9D16: data_out = 8'h87;
                    16'h9D17: data_out = 8'h86;
                    16'h9D18: data_out = 8'h85;
                    16'h9D19: data_out = 8'h84;
                    16'h9D1A: data_out = 8'h83;
                    16'h9D1B: data_out = 8'h82;
                    16'h9D1C: data_out = 8'h81;
                    16'h9D1D: data_out = 8'h0;
                    16'h9D1E: data_out = 8'h1;
                    16'h9D1F: data_out = 8'h2;
                    16'h9D20: data_out = 8'h3;
                    16'h9D21: data_out = 8'h4;
                    16'h9D22: data_out = 8'h5;
                    16'h9D23: data_out = 8'h6;
                    16'h9D24: data_out = 8'h7;
                    16'h9D25: data_out = 8'h8;
                    16'h9D26: data_out = 8'h9;
                    16'h9D27: data_out = 8'hA;
                    16'h9D28: data_out = 8'hB;
                    16'h9D29: data_out = 8'hC;
                    16'h9D2A: data_out = 8'hD;
                    16'h9D2B: data_out = 8'hE;
                    16'h9D2C: data_out = 8'hF;
                    16'h9D2D: data_out = 8'h10;
                    16'h9D2E: data_out = 8'h11;
                    16'h9D2F: data_out = 8'h12;
                    16'h9D30: data_out = 8'h13;
                    16'h9D31: data_out = 8'h14;
                    16'h9D32: data_out = 8'h15;
                    16'h9D33: data_out = 8'h16;
                    16'h9D34: data_out = 8'h17;
                    16'h9D35: data_out = 8'h18;
                    16'h9D36: data_out = 8'h19;
                    16'h9D37: data_out = 8'h1A;
                    16'h9D38: data_out = 8'h1B;
                    16'h9D39: data_out = 8'h1C;
                    16'h9D3A: data_out = 8'h1D;
                    16'h9D3B: data_out = 8'h1E;
                    16'h9D3C: data_out = 8'h1F;
                    16'h9D3D: data_out = 8'h20;
                    16'h9D3E: data_out = 8'h21;
                    16'h9D3F: data_out = 8'h22;
                    16'h9D40: data_out = 8'h23;
                    16'h9D41: data_out = 8'h24;
                    16'h9D42: data_out = 8'h25;
                    16'h9D43: data_out = 8'h26;
                    16'h9D44: data_out = 8'h27;
                    16'h9D45: data_out = 8'h28;
                    16'h9D46: data_out = 8'h29;
                    16'h9D47: data_out = 8'h2A;
                    16'h9D48: data_out = 8'h2B;
                    16'h9D49: data_out = 8'h2C;
                    16'h9D4A: data_out = 8'h2D;
                    16'h9D4B: data_out = 8'h2E;
                    16'h9D4C: data_out = 8'h2F;
                    16'h9D4D: data_out = 8'h30;
                    16'h9D4E: data_out = 8'h31;
                    16'h9D4F: data_out = 8'h32;
                    16'h9D50: data_out = 8'h33;
                    16'h9D51: data_out = 8'h34;
                    16'h9D52: data_out = 8'h35;
                    16'h9D53: data_out = 8'h36;
                    16'h9D54: data_out = 8'h37;
                    16'h9D55: data_out = 8'h38;
                    16'h9D56: data_out = 8'h39;
                    16'h9D57: data_out = 8'h3A;
                    16'h9D58: data_out = 8'h3B;
                    16'h9D59: data_out = 8'h3C;
                    16'h9D5A: data_out = 8'h3D;
                    16'h9D5B: data_out = 8'h3E;
                    16'h9D5C: data_out = 8'h3F;
                    16'h9D5D: data_out = 8'h40;
                    16'h9D5E: data_out = 8'h41;
                    16'h9D5F: data_out = 8'h42;
                    16'h9D60: data_out = 8'h43;
                    16'h9D61: data_out = 8'h44;
                    16'h9D62: data_out = 8'h45;
                    16'h9D63: data_out = 8'h46;
                    16'h9D64: data_out = 8'h47;
                    16'h9D65: data_out = 8'h48;
                    16'h9D66: data_out = 8'h49;
                    16'h9D67: data_out = 8'h4A;
                    16'h9D68: data_out = 8'h4B;
                    16'h9D69: data_out = 8'h4C;
                    16'h9D6A: data_out = 8'h4D;
                    16'h9D6B: data_out = 8'h4E;
                    16'h9D6C: data_out = 8'h4F;
                    16'h9D6D: data_out = 8'h50;
                    16'h9D6E: data_out = 8'h51;
                    16'h9D6F: data_out = 8'h52;
                    16'h9D70: data_out = 8'h53;
                    16'h9D71: data_out = 8'h54;
                    16'h9D72: data_out = 8'h55;
                    16'h9D73: data_out = 8'h56;
                    16'h9D74: data_out = 8'h57;
                    16'h9D75: data_out = 8'h58;
                    16'h9D76: data_out = 8'h59;
                    16'h9D77: data_out = 8'h5A;
                    16'h9D78: data_out = 8'h5B;
                    16'h9D79: data_out = 8'h5C;
                    16'h9D7A: data_out = 8'h5D;
                    16'h9D7B: data_out = 8'h5E;
                    16'h9D7C: data_out = 8'h5F;
                    16'h9D7D: data_out = 8'h60;
                    16'h9D7E: data_out = 8'h61;
                    16'h9D7F: data_out = 8'h62;
                    16'h9D80: data_out = 8'h9D;
                    16'h9D81: data_out = 8'h9E;
                    16'h9D82: data_out = 8'h9F;
                    16'h9D83: data_out = 8'hA0;
                    16'h9D84: data_out = 8'hA1;
                    16'h9D85: data_out = 8'hA2;
                    16'h9D86: data_out = 8'hA3;
                    16'h9D87: data_out = 8'hA4;
                    16'h9D88: data_out = 8'hA5;
                    16'h9D89: data_out = 8'hA6;
                    16'h9D8A: data_out = 8'hA7;
                    16'h9D8B: data_out = 8'hA8;
                    16'h9D8C: data_out = 8'hA9;
                    16'h9D8D: data_out = 8'hAA;
                    16'h9D8E: data_out = 8'hAB;
                    16'h9D8F: data_out = 8'hAC;
                    16'h9D90: data_out = 8'hAD;
                    16'h9D91: data_out = 8'hAE;
                    16'h9D92: data_out = 8'hAF;
                    16'h9D93: data_out = 8'hB0;
                    16'h9D94: data_out = 8'hB1;
                    16'h9D95: data_out = 8'hB2;
                    16'h9D96: data_out = 8'hB3;
                    16'h9D97: data_out = 8'hB4;
                    16'h9D98: data_out = 8'hB5;
                    16'h9D99: data_out = 8'hB6;
                    16'h9D9A: data_out = 8'hB7;
                    16'h9D9B: data_out = 8'hB8;
                    16'h9D9C: data_out = 8'hB9;
                    16'h9D9D: data_out = 8'hBA;
                    16'h9D9E: data_out = 8'hBB;
                    16'h9D9F: data_out = 8'hBC;
                    16'h9DA0: data_out = 8'hBD;
                    16'h9DA1: data_out = 8'hBE;
                    16'h9DA2: data_out = 8'hBF;
                    16'h9DA3: data_out = 8'hC0;
                    16'h9DA4: data_out = 8'hC1;
                    16'h9DA5: data_out = 8'hC2;
                    16'h9DA6: data_out = 8'hC3;
                    16'h9DA7: data_out = 8'hC4;
                    16'h9DA8: data_out = 8'hC5;
                    16'h9DA9: data_out = 8'hC6;
                    16'h9DAA: data_out = 8'hC7;
                    16'h9DAB: data_out = 8'hC8;
                    16'h9DAC: data_out = 8'hC9;
                    16'h9DAD: data_out = 8'hCA;
                    16'h9DAE: data_out = 8'hCB;
                    16'h9DAF: data_out = 8'hCC;
                    16'h9DB0: data_out = 8'hCD;
                    16'h9DB1: data_out = 8'hCE;
                    16'h9DB2: data_out = 8'hCF;
                    16'h9DB3: data_out = 8'hD0;
                    16'h9DB4: data_out = 8'hD1;
                    16'h9DB5: data_out = 8'hD2;
                    16'h9DB6: data_out = 8'hD3;
                    16'h9DB7: data_out = 8'hD4;
                    16'h9DB8: data_out = 8'hD5;
                    16'h9DB9: data_out = 8'hD6;
                    16'h9DBA: data_out = 8'hD7;
                    16'h9DBB: data_out = 8'hD8;
                    16'h9DBC: data_out = 8'hD9;
                    16'h9DBD: data_out = 8'hDA;
                    16'h9DBE: data_out = 8'hDB;
                    16'h9DBF: data_out = 8'hDC;
                    16'h9DC0: data_out = 8'hDD;
                    16'h9DC1: data_out = 8'hDE;
                    16'h9DC2: data_out = 8'hDF;
                    16'h9DC3: data_out = 8'hE0;
                    16'h9DC4: data_out = 8'hE1;
                    16'h9DC5: data_out = 8'hE2;
                    16'h9DC6: data_out = 8'hE3;
                    16'h9DC7: data_out = 8'hE4;
                    16'h9DC8: data_out = 8'hE5;
                    16'h9DC9: data_out = 8'hE6;
                    16'h9DCA: data_out = 8'hE7;
                    16'h9DCB: data_out = 8'hE8;
                    16'h9DCC: data_out = 8'hE9;
                    16'h9DCD: data_out = 8'hEA;
                    16'h9DCE: data_out = 8'hEB;
                    16'h9DCF: data_out = 8'hEC;
                    16'h9DD0: data_out = 8'hED;
                    16'h9DD1: data_out = 8'hEE;
                    16'h9DD2: data_out = 8'hEF;
                    16'h9DD3: data_out = 8'hF0;
                    16'h9DD4: data_out = 8'hF1;
                    16'h9DD5: data_out = 8'hF2;
                    16'h9DD6: data_out = 8'hF3;
                    16'h9DD7: data_out = 8'hF4;
                    16'h9DD8: data_out = 8'hF5;
                    16'h9DD9: data_out = 8'hF6;
                    16'h9DDA: data_out = 8'hF7;
                    16'h9DDB: data_out = 8'hF8;
                    16'h9DDC: data_out = 8'hF9;
                    16'h9DDD: data_out = 8'hFA;
                    16'h9DDE: data_out = 8'hFB;
                    16'h9DDF: data_out = 8'hFC;
                    16'h9DE0: data_out = 8'hFD;
                    16'h9DE1: data_out = 8'hFE;
                    16'h9DE2: data_out = 8'hFF;
                    16'h9DE3: data_out = 8'h80;
                    16'h9DE4: data_out = 8'h81;
                    16'h9DE5: data_out = 8'h82;
                    16'h9DE6: data_out = 8'h83;
                    16'h9DE7: data_out = 8'h84;
                    16'h9DE8: data_out = 8'h85;
                    16'h9DE9: data_out = 8'h86;
                    16'h9DEA: data_out = 8'h87;
                    16'h9DEB: data_out = 8'h88;
                    16'h9DEC: data_out = 8'h89;
                    16'h9DED: data_out = 8'h8A;
                    16'h9DEE: data_out = 8'h8B;
                    16'h9DEF: data_out = 8'h8C;
                    16'h9DF0: data_out = 8'h8D;
                    16'h9DF1: data_out = 8'h8E;
                    16'h9DF2: data_out = 8'h8F;
                    16'h9DF3: data_out = 8'h90;
                    16'h9DF4: data_out = 8'h91;
                    16'h9DF5: data_out = 8'h92;
                    16'h9DF6: data_out = 8'h93;
                    16'h9DF7: data_out = 8'h94;
                    16'h9DF8: data_out = 8'h95;
                    16'h9DF9: data_out = 8'h96;
                    16'h9DFA: data_out = 8'h97;
                    16'h9DFB: data_out = 8'h98;
                    16'h9DFC: data_out = 8'h99;
                    16'h9DFD: data_out = 8'h9A;
                    16'h9DFE: data_out = 8'h9B;
                    16'h9DFF: data_out = 8'h9C;
                    16'h9E00: data_out = 8'h9E;
                    16'h9E01: data_out = 8'h9D;
                    16'h9E02: data_out = 8'h9C;
                    16'h9E03: data_out = 8'h9B;
                    16'h9E04: data_out = 8'h9A;
                    16'h9E05: data_out = 8'h99;
                    16'h9E06: data_out = 8'h98;
                    16'h9E07: data_out = 8'h97;
                    16'h9E08: data_out = 8'h96;
                    16'h9E09: data_out = 8'h95;
                    16'h9E0A: data_out = 8'h94;
                    16'h9E0B: data_out = 8'h93;
                    16'h9E0C: data_out = 8'h92;
                    16'h9E0D: data_out = 8'h91;
                    16'h9E0E: data_out = 8'h90;
                    16'h9E0F: data_out = 8'h8F;
                    16'h9E10: data_out = 8'h8E;
                    16'h9E11: data_out = 8'h8D;
                    16'h9E12: data_out = 8'h8C;
                    16'h9E13: data_out = 8'h8B;
                    16'h9E14: data_out = 8'h8A;
                    16'h9E15: data_out = 8'h89;
                    16'h9E16: data_out = 8'h88;
                    16'h9E17: data_out = 8'h87;
                    16'h9E18: data_out = 8'h86;
                    16'h9E19: data_out = 8'h85;
                    16'h9E1A: data_out = 8'h84;
                    16'h9E1B: data_out = 8'h83;
                    16'h9E1C: data_out = 8'h82;
                    16'h9E1D: data_out = 8'h81;
                    16'h9E1E: data_out = 8'h0;
                    16'h9E1F: data_out = 8'h1;
                    16'h9E20: data_out = 8'h2;
                    16'h9E21: data_out = 8'h3;
                    16'h9E22: data_out = 8'h4;
                    16'h9E23: data_out = 8'h5;
                    16'h9E24: data_out = 8'h6;
                    16'h9E25: data_out = 8'h7;
                    16'h9E26: data_out = 8'h8;
                    16'h9E27: data_out = 8'h9;
                    16'h9E28: data_out = 8'hA;
                    16'h9E29: data_out = 8'hB;
                    16'h9E2A: data_out = 8'hC;
                    16'h9E2B: data_out = 8'hD;
                    16'h9E2C: data_out = 8'hE;
                    16'h9E2D: data_out = 8'hF;
                    16'h9E2E: data_out = 8'h10;
                    16'h9E2F: data_out = 8'h11;
                    16'h9E30: data_out = 8'h12;
                    16'h9E31: data_out = 8'h13;
                    16'h9E32: data_out = 8'h14;
                    16'h9E33: data_out = 8'h15;
                    16'h9E34: data_out = 8'h16;
                    16'h9E35: data_out = 8'h17;
                    16'h9E36: data_out = 8'h18;
                    16'h9E37: data_out = 8'h19;
                    16'h9E38: data_out = 8'h1A;
                    16'h9E39: data_out = 8'h1B;
                    16'h9E3A: data_out = 8'h1C;
                    16'h9E3B: data_out = 8'h1D;
                    16'h9E3C: data_out = 8'h1E;
                    16'h9E3D: data_out = 8'h1F;
                    16'h9E3E: data_out = 8'h20;
                    16'h9E3F: data_out = 8'h21;
                    16'h9E40: data_out = 8'h22;
                    16'h9E41: data_out = 8'h23;
                    16'h9E42: data_out = 8'h24;
                    16'h9E43: data_out = 8'h25;
                    16'h9E44: data_out = 8'h26;
                    16'h9E45: data_out = 8'h27;
                    16'h9E46: data_out = 8'h28;
                    16'h9E47: data_out = 8'h29;
                    16'h9E48: data_out = 8'h2A;
                    16'h9E49: data_out = 8'h2B;
                    16'h9E4A: data_out = 8'h2C;
                    16'h9E4B: data_out = 8'h2D;
                    16'h9E4C: data_out = 8'h2E;
                    16'h9E4D: data_out = 8'h2F;
                    16'h9E4E: data_out = 8'h30;
                    16'h9E4F: data_out = 8'h31;
                    16'h9E50: data_out = 8'h32;
                    16'h9E51: data_out = 8'h33;
                    16'h9E52: data_out = 8'h34;
                    16'h9E53: data_out = 8'h35;
                    16'h9E54: data_out = 8'h36;
                    16'h9E55: data_out = 8'h37;
                    16'h9E56: data_out = 8'h38;
                    16'h9E57: data_out = 8'h39;
                    16'h9E58: data_out = 8'h3A;
                    16'h9E59: data_out = 8'h3B;
                    16'h9E5A: data_out = 8'h3C;
                    16'h9E5B: data_out = 8'h3D;
                    16'h9E5C: data_out = 8'h3E;
                    16'h9E5D: data_out = 8'h3F;
                    16'h9E5E: data_out = 8'h40;
                    16'h9E5F: data_out = 8'h41;
                    16'h9E60: data_out = 8'h42;
                    16'h9E61: data_out = 8'h43;
                    16'h9E62: data_out = 8'h44;
                    16'h9E63: data_out = 8'h45;
                    16'h9E64: data_out = 8'h46;
                    16'h9E65: data_out = 8'h47;
                    16'h9E66: data_out = 8'h48;
                    16'h9E67: data_out = 8'h49;
                    16'h9E68: data_out = 8'h4A;
                    16'h9E69: data_out = 8'h4B;
                    16'h9E6A: data_out = 8'h4C;
                    16'h9E6B: data_out = 8'h4D;
                    16'h9E6C: data_out = 8'h4E;
                    16'h9E6D: data_out = 8'h4F;
                    16'h9E6E: data_out = 8'h50;
                    16'h9E6F: data_out = 8'h51;
                    16'h9E70: data_out = 8'h52;
                    16'h9E71: data_out = 8'h53;
                    16'h9E72: data_out = 8'h54;
                    16'h9E73: data_out = 8'h55;
                    16'h9E74: data_out = 8'h56;
                    16'h9E75: data_out = 8'h57;
                    16'h9E76: data_out = 8'h58;
                    16'h9E77: data_out = 8'h59;
                    16'h9E78: data_out = 8'h5A;
                    16'h9E79: data_out = 8'h5B;
                    16'h9E7A: data_out = 8'h5C;
                    16'h9E7B: data_out = 8'h5D;
                    16'h9E7C: data_out = 8'h5E;
                    16'h9E7D: data_out = 8'h5F;
                    16'h9E7E: data_out = 8'h60;
                    16'h9E7F: data_out = 8'h61;
                    16'h9E80: data_out = 8'h9E;
                    16'h9E81: data_out = 8'h9F;
                    16'h9E82: data_out = 8'hA0;
                    16'h9E83: data_out = 8'hA1;
                    16'h9E84: data_out = 8'hA2;
                    16'h9E85: data_out = 8'hA3;
                    16'h9E86: data_out = 8'hA4;
                    16'h9E87: data_out = 8'hA5;
                    16'h9E88: data_out = 8'hA6;
                    16'h9E89: data_out = 8'hA7;
                    16'h9E8A: data_out = 8'hA8;
                    16'h9E8B: data_out = 8'hA9;
                    16'h9E8C: data_out = 8'hAA;
                    16'h9E8D: data_out = 8'hAB;
                    16'h9E8E: data_out = 8'hAC;
                    16'h9E8F: data_out = 8'hAD;
                    16'h9E90: data_out = 8'hAE;
                    16'h9E91: data_out = 8'hAF;
                    16'h9E92: data_out = 8'hB0;
                    16'h9E93: data_out = 8'hB1;
                    16'h9E94: data_out = 8'hB2;
                    16'h9E95: data_out = 8'hB3;
                    16'h9E96: data_out = 8'hB4;
                    16'h9E97: data_out = 8'hB5;
                    16'h9E98: data_out = 8'hB6;
                    16'h9E99: data_out = 8'hB7;
                    16'h9E9A: data_out = 8'hB8;
                    16'h9E9B: data_out = 8'hB9;
                    16'h9E9C: data_out = 8'hBA;
                    16'h9E9D: data_out = 8'hBB;
                    16'h9E9E: data_out = 8'hBC;
                    16'h9E9F: data_out = 8'hBD;
                    16'h9EA0: data_out = 8'hBE;
                    16'h9EA1: data_out = 8'hBF;
                    16'h9EA2: data_out = 8'hC0;
                    16'h9EA3: data_out = 8'hC1;
                    16'h9EA4: data_out = 8'hC2;
                    16'h9EA5: data_out = 8'hC3;
                    16'h9EA6: data_out = 8'hC4;
                    16'h9EA7: data_out = 8'hC5;
                    16'h9EA8: data_out = 8'hC6;
                    16'h9EA9: data_out = 8'hC7;
                    16'h9EAA: data_out = 8'hC8;
                    16'h9EAB: data_out = 8'hC9;
                    16'h9EAC: data_out = 8'hCA;
                    16'h9EAD: data_out = 8'hCB;
                    16'h9EAE: data_out = 8'hCC;
                    16'h9EAF: data_out = 8'hCD;
                    16'h9EB0: data_out = 8'hCE;
                    16'h9EB1: data_out = 8'hCF;
                    16'h9EB2: data_out = 8'hD0;
                    16'h9EB3: data_out = 8'hD1;
                    16'h9EB4: data_out = 8'hD2;
                    16'h9EB5: data_out = 8'hD3;
                    16'h9EB6: data_out = 8'hD4;
                    16'h9EB7: data_out = 8'hD5;
                    16'h9EB8: data_out = 8'hD6;
                    16'h9EB9: data_out = 8'hD7;
                    16'h9EBA: data_out = 8'hD8;
                    16'h9EBB: data_out = 8'hD9;
                    16'h9EBC: data_out = 8'hDA;
                    16'h9EBD: data_out = 8'hDB;
                    16'h9EBE: data_out = 8'hDC;
                    16'h9EBF: data_out = 8'hDD;
                    16'h9EC0: data_out = 8'hDE;
                    16'h9EC1: data_out = 8'hDF;
                    16'h9EC2: data_out = 8'hE0;
                    16'h9EC3: data_out = 8'hE1;
                    16'h9EC4: data_out = 8'hE2;
                    16'h9EC5: data_out = 8'hE3;
                    16'h9EC6: data_out = 8'hE4;
                    16'h9EC7: data_out = 8'hE5;
                    16'h9EC8: data_out = 8'hE6;
                    16'h9EC9: data_out = 8'hE7;
                    16'h9ECA: data_out = 8'hE8;
                    16'h9ECB: data_out = 8'hE9;
                    16'h9ECC: data_out = 8'hEA;
                    16'h9ECD: data_out = 8'hEB;
                    16'h9ECE: data_out = 8'hEC;
                    16'h9ECF: data_out = 8'hED;
                    16'h9ED0: data_out = 8'hEE;
                    16'h9ED1: data_out = 8'hEF;
                    16'h9ED2: data_out = 8'hF0;
                    16'h9ED3: data_out = 8'hF1;
                    16'h9ED4: data_out = 8'hF2;
                    16'h9ED5: data_out = 8'hF3;
                    16'h9ED6: data_out = 8'hF4;
                    16'h9ED7: data_out = 8'hF5;
                    16'h9ED8: data_out = 8'hF6;
                    16'h9ED9: data_out = 8'hF7;
                    16'h9EDA: data_out = 8'hF8;
                    16'h9EDB: data_out = 8'hF9;
                    16'h9EDC: data_out = 8'hFA;
                    16'h9EDD: data_out = 8'hFB;
                    16'h9EDE: data_out = 8'hFC;
                    16'h9EDF: data_out = 8'hFD;
                    16'h9EE0: data_out = 8'hFE;
                    16'h9EE1: data_out = 8'hFF;
                    16'h9EE2: data_out = 8'h80;
                    16'h9EE3: data_out = 8'h81;
                    16'h9EE4: data_out = 8'h82;
                    16'h9EE5: data_out = 8'h83;
                    16'h9EE6: data_out = 8'h84;
                    16'h9EE7: data_out = 8'h85;
                    16'h9EE8: data_out = 8'h86;
                    16'h9EE9: data_out = 8'h87;
                    16'h9EEA: data_out = 8'h88;
                    16'h9EEB: data_out = 8'h89;
                    16'h9EEC: data_out = 8'h8A;
                    16'h9EED: data_out = 8'h8B;
                    16'h9EEE: data_out = 8'h8C;
                    16'h9EEF: data_out = 8'h8D;
                    16'h9EF0: data_out = 8'h8E;
                    16'h9EF1: data_out = 8'h8F;
                    16'h9EF2: data_out = 8'h90;
                    16'h9EF3: data_out = 8'h91;
                    16'h9EF4: data_out = 8'h92;
                    16'h9EF5: data_out = 8'h93;
                    16'h9EF6: data_out = 8'h94;
                    16'h9EF7: data_out = 8'h95;
                    16'h9EF8: data_out = 8'h96;
                    16'h9EF9: data_out = 8'h97;
                    16'h9EFA: data_out = 8'h98;
                    16'h9EFB: data_out = 8'h99;
                    16'h9EFC: data_out = 8'h9A;
                    16'h9EFD: data_out = 8'h9B;
                    16'h9EFE: data_out = 8'h9C;
                    16'h9EFF: data_out = 8'h9D;
                    16'h9F00: data_out = 8'h9F;
                    16'h9F01: data_out = 8'h9E;
                    16'h9F02: data_out = 8'h9D;
                    16'h9F03: data_out = 8'h9C;
                    16'h9F04: data_out = 8'h9B;
                    16'h9F05: data_out = 8'h9A;
                    16'h9F06: data_out = 8'h99;
                    16'h9F07: data_out = 8'h98;
                    16'h9F08: data_out = 8'h97;
                    16'h9F09: data_out = 8'h96;
                    16'h9F0A: data_out = 8'h95;
                    16'h9F0B: data_out = 8'h94;
                    16'h9F0C: data_out = 8'h93;
                    16'h9F0D: data_out = 8'h92;
                    16'h9F0E: data_out = 8'h91;
                    16'h9F0F: data_out = 8'h90;
                    16'h9F10: data_out = 8'h8F;
                    16'h9F11: data_out = 8'h8E;
                    16'h9F12: data_out = 8'h8D;
                    16'h9F13: data_out = 8'h8C;
                    16'h9F14: data_out = 8'h8B;
                    16'h9F15: data_out = 8'h8A;
                    16'h9F16: data_out = 8'h89;
                    16'h9F17: data_out = 8'h88;
                    16'h9F18: data_out = 8'h87;
                    16'h9F19: data_out = 8'h86;
                    16'h9F1A: data_out = 8'h85;
                    16'h9F1B: data_out = 8'h84;
                    16'h9F1C: data_out = 8'h83;
                    16'h9F1D: data_out = 8'h82;
                    16'h9F1E: data_out = 8'h81;
                    16'h9F1F: data_out = 8'h0;
                    16'h9F20: data_out = 8'h1;
                    16'h9F21: data_out = 8'h2;
                    16'h9F22: data_out = 8'h3;
                    16'h9F23: data_out = 8'h4;
                    16'h9F24: data_out = 8'h5;
                    16'h9F25: data_out = 8'h6;
                    16'h9F26: data_out = 8'h7;
                    16'h9F27: data_out = 8'h8;
                    16'h9F28: data_out = 8'h9;
                    16'h9F29: data_out = 8'hA;
                    16'h9F2A: data_out = 8'hB;
                    16'h9F2B: data_out = 8'hC;
                    16'h9F2C: data_out = 8'hD;
                    16'h9F2D: data_out = 8'hE;
                    16'h9F2E: data_out = 8'hF;
                    16'h9F2F: data_out = 8'h10;
                    16'h9F30: data_out = 8'h11;
                    16'h9F31: data_out = 8'h12;
                    16'h9F32: data_out = 8'h13;
                    16'h9F33: data_out = 8'h14;
                    16'h9F34: data_out = 8'h15;
                    16'h9F35: data_out = 8'h16;
                    16'h9F36: data_out = 8'h17;
                    16'h9F37: data_out = 8'h18;
                    16'h9F38: data_out = 8'h19;
                    16'h9F39: data_out = 8'h1A;
                    16'h9F3A: data_out = 8'h1B;
                    16'h9F3B: data_out = 8'h1C;
                    16'h9F3C: data_out = 8'h1D;
                    16'h9F3D: data_out = 8'h1E;
                    16'h9F3E: data_out = 8'h1F;
                    16'h9F3F: data_out = 8'h20;
                    16'h9F40: data_out = 8'h21;
                    16'h9F41: data_out = 8'h22;
                    16'h9F42: data_out = 8'h23;
                    16'h9F43: data_out = 8'h24;
                    16'h9F44: data_out = 8'h25;
                    16'h9F45: data_out = 8'h26;
                    16'h9F46: data_out = 8'h27;
                    16'h9F47: data_out = 8'h28;
                    16'h9F48: data_out = 8'h29;
                    16'h9F49: data_out = 8'h2A;
                    16'h9F4A: data_out = 8'h2B;
                    16'h9F4B: data_out = 8'h2C;
                    16'h9F4C: data_out = 8'h2D;
                    16'h9F4D: data_out = 8'h2E;
                    16'h9F4E: data_out = 8'h2F;
                    16'h9F4F: data_out = 8'h30;
                    16'h9F50: data_out = 8'h31;
                    16'h9F51: data_out = 8'h32;
                    16'h9F52: data_out = 8'h33;
                    16'h9F53: data_out = 8'h34;
                    16'h9F54: data_out = 8'h35;
                    16'h9F55: data_out = 8'h36;
                    16'h9F56: data_out = 8'h37;
                    16'h9F57: data_out = 8'h38;
                    16'h9F58: data_out = 8'h39;
                    16'h9F59: data_out = 8'h3A;
                    16'h9F5A: data_out = 8'h3B;
                    16'h9F5B: data_out = 8'h3C;
                    16'h9F5C: data_out = 8'h3D;
                    16'h9F5D: data_out = 8'h3E;
                    16'h9F5E: data_out = 8'h3F;
                    16'h9F5F: data_out = 8'h40;
                    16'h9F60: data_out = 8'h41;
                    16'h9F61: data_out = 8'h42;
                    16'h9F62: data_out = 8'h43;
                    16'h9F63: data_out = 8'h44;
                    16'h9F64: data_out = 8'h45;
                    16'h9F65: data_out = 8'h46;
                    16'h9F66: data_out = 8'h47;
                    16'h9F67: data_out = 8'h48;
                    16'h9F68: data_out = 8'h49;
                    16'h9F69: data_out = 8'h4A;
                    16'h9F6A: data_out = 8'h4B;
                    16'h9F6B: data_out = 8'h4C;
                    16'h9F6C: data_out = 8'h4D;
                    16'h9F6D: data_out = 8'h4E;
                    16'h9F6E: data_out = 8'h4F;
                    16'h9F6F: data_out = 8'h50;
                    16'h9F70: data_out = 8'h51;
                    16'h9F71: data_out = 8'h52;
                    16'h9F72: data_out = 8'h53;
                    16'h9F73: data_out = 8'h54;
                    16'h9F74: data_out = 8'h55;
                    16'h9F75: data_out = 8'h56;
                    16'h9F76: data_out = 8'h57;
                    16'h9F77: data_out = 8'h58;
                    16'h9F78: data_out = 8'h59;
                    16'h9F79: data_out = 8'h5A;
                    16'h9F7A: data_out = 8'h5B;
                    16'h9F7B: data_out = 8'h5C;
                    16'h9F7C: data_out = 8'h5D;
                    16'h9F7D: data_out = 8'h5E;
                    16'h9F7E: data_out = 8'h5F;
                    16'h9F7F: data_out = 8'h60;
                    16'h9F80: data_out = 8'h9F;
                    16'h9F81: data_out = 8'hA0;
                    16'h9F82: data_out = 8'hA1;
                    16'h9F83: data_out = 8'hA2;
                    16'h9F84: data_out = 8'hA3;
                    16'h9F85: data_out = 8'hA4;
                    16'h9F86: data_out = 8'hA5;
                    16'h9F87: data_out = 8'hA6;
                    16'h9F88: data_out = 8'hA7;
                    16'h9F89: data_out = 8'hA8;
                    16'h9F8A: data_out = 8'hA9;
                    16'h9F8B: data_out = 8'hAA;
                    16'h9F8C: data_out = 8'hAB;
                    16'h9F8D: data_out = 8'hAC;
                    16'h9F8E: data_out = 8'hAD;
                    16'h9F8F: data_out = 8'hAE;
                    16'h9F90: data_out = 8'hAF;
                    16'h9F91: data_out = 8'hB0;
                    16'h9F92: data_out = 8'hB1;
                    16'h9F93: data_out = 8'hB2;
                    16'h9F94: data_out = 8'hB3;
                    16'h9F95: data_out = 8'hB4;
                    16'h9F96: data_out = 8'hB5;
                    16'h9F97: data_out = 8'hB6;
                    16'h9F98: data_out = 8'hB7;
                    16'h9F99: data_out = 8'hB8;
                    16'h9F9A: data_out = 8'hB9;
                    16'h9F9B: data_out = 8'hBA;
                    16'h9F9C: data_out = 8'hBB;
                    16'h9F9D: data_out = 8'hBC;
                    16'h9F9E: data_out = 8'hBD;
                    16'h9F9F: data_out = 8'hBE;
                    16'h9FA0: data_out = 8'hBF;
                    16'h9FA1: data_out = 8'hC0;
                    16'h9FA2: data_out = 8'hC1;
                    16'h9FA3: data_out = 8'hC2;
                    16'h9FA4: data_out = 8'hC3;
                    16'h9FA5: data_out = 8'hC4;
                    16'h9FA6: data_out = 8'hC5;
                    16'h9FA7: data_out = 8'hC6;
                    16'h9FA8: data_out = 8'hC7;
                    16'h9FA9: data_out = 8'hC8;
                    16'h9FAA: data_out = 8'hC9;
                    16'h9FAB: data_out = 8'hCA;
                    16'h9FAC: data_out = 8'hCB;
                    16'h9FAD: data_out = 8'hCC;
                    16'h9FAE: data_out = 8'hCD;
                    16'h9FAF: data_out = 8'hCE;
                    16'h9FB0: data_out = 8'hCF;
                    16'h9FB1: data_out = 8'hD0;
                    16'h9FB2: data_out = 8'hD1;
                    16'h9FB3: data_out = 8'hD2;
                    16'h9FB4: data_out = 8'hD3;
                    16'h9FB5: data_out = 8'hD4;
                    16'h9FB6: data_out = 8'hD5;
                    16'h9FB7: data_out = 8'hD6;
                    16'h9FB8: data_out = 8'hD7;
                    16'h9FB9: data_out = 8'hD8;
                    16'h9FBA: data_out = 8'hD9;
                    16'h9FBB: data_out = 8'hDA;
                    16'h9FBC: data_out = 8'hDB;
                    16'h9FBD: data_out = 8'hDC;
                    16'h9FBE: data_out = 8'hDD;
                    16'h9FBF: data_out = 8'hDE;
                    16'h9FC0: data_out = 8'hDF;
                    16'h9FC1: data_out = 8'hE0;
                    16'h9FC2: data_out = 8'hE1;
                    16'h9FC3: data_out = 8'hE2;
                    16'h9FC4: data_out = 8'hE3;
                    16'h9FC5: data_out = 8'hE4;
                    16'h9FC6: data_out = 8'hE5;
                    16'h9FC7: data_out = 8'hE6;
                    16'h9FC8: data_out = 8'hE7;
                    16'h9FC9: data_out = 8'hE8;
                    16'h9FCA: data_out = 8'hE9;
                    16'h9FCB: data_out = 8'hEA;
                    16'h9FCC: data_out = 8'hEB;
                    16'h9FCD: data_out = 8'hEC;
                    16'h9FCE: data_out = 8'hED;
                    16'h9FCF: data_out = 8'hEE;
                    16'h9FD0: data_out = 8'hEF;
                    16'h9FD1: data_out = 8'hF0;
                    16'h9FD2: data_out = 8'hF1;
                    16'h9FD3: data_out = 8'hF2;
                    16'h9FD4: data_out = 8'hF3;
                    16'h9FD5: data_out = 8'hF4;
                    16'h9FD6: data_out = 8'hF5;
                    16'h9FD7: data_out = 8'hF6;
                    16'h9FD8: data_out = 8'hF7;
                    16'h9FD9: data_out = 8'hF8;
                    16'h9FDA: data_out = 8'hF9;
                    16'h9FDB: data_out = 8'hFA;
                    16'h9FDC: data_out = 8'hFB;
                    16'h9FDD: data_out = 8'hFC;
                    16'h9FDE: data_out = 8'hFD;
                    16'h9FDF: data_out = 8'hFE;
                    16'h9FE0: data_out = 8'hFF;
                    16'h9FE1: data_out = 8'h80;
                    16'h9FE2: data_out = 8'h81;
                    16'h9FE3: data_out = 8'h82;
                    16'h9FE4: data_out = 8'h83;
                    16'h9FE5: data_out = 8'h84;
                    16'h9FE6: data_out = 8'h85;
                    16'h9FE7: data_out = 8'h86;
                    16'h9FE8: data_out = 8'h87;
                    16'h9FE9: data_out = 8'h88;
                    16'h9FEA: data_out = 8'h89;
                    16'h9FEB: data_out = 8'h8A;
                    16'h9FEC: data_out = 8'h8B;
                    16'h9FED: data_out = 8'h8C;
                    16'h9FEE: data_out = 8'h8D;
                    16'h9FEF: data_out = 8'h8E;
                    16'h9FF0: data_out = 8'h8F;
                    16'h9FF1: data_out = 8'h90;
                    16'h9FF2: data_out = 8'h91;
                    16'h9FF3: data_out = 8'h92;
                    16'h9FF4: data_out = 8'h93;
                    16'h9FF5: data_out = 8'h94;
                    16'h9FF6: data_out = 8'h95;
                    16'h9FF7: data_out = 8'h96;
                    16'h9FF8: data_out = 8'h97;
                    16'h9FF9: data_out = 8'h98;
                    16'h9FFA: data_out = 8'h99;
                    16'h9FFB: data_out = 8'h9A;
                    16'h9FFC: data_out = 8'h9B;
                    16'h9FFD: data_out = 8'h9C;
                    16'h9FFE: data_out = 8'h9D;
                    16'h9FFF: data_out = 8'h9E;
                    16'hA000: data_out = 8'hA0;
                    16'hA001: data_out = 8'h9F;
                    16'hA002: data_out = 8'h9E;
                    16'hA003: data_out = 8'h9D;
                    16'hA004: data_out = 8'h9C;
                    16'hA005: data_out = 8'h9B;
                    16'hA006: data_out = 8'h9A;
                    16'hA007: data_out = 8'h99;
                    16'hA008: data_out = 8'h98;
                    16'hA009: data_out = 8'h97;
                    16'hA00A: data_out = 8'h96;
                    16'hA00B: data_out = 8'h95;
                    16'hA00C: data_out = 8'h94;
                    16'hA00D: data_out = 8'h93;
                    16'hA00E: data_out = 8'h92;
                    16'hA00F: data_out = 8'h91;
                    16'hA010: data_out = 8'h90;
                    16'hA011: data_out = 8'h8F;
                    16'hA012: data_out = 8'h8E;
                    16'hA013: data_out = 8'h8D;
                    16'hA014: data_out = 8'h8C;
                    16'hA015: data_out = 8'h8B;
                    16'hA016: data_out = 8'h8A;
                    16'hA017: data_out = 8'h89;
                    16'hA018: data_out = 8'h88;
                    16'hA019: data_out = 8'h87;
                    16'hA01A: data_out = 8'h86;
                    16'hA01B: data_out = 8'h85;
                    16'hA01C: data_out = 8'h84;
                    16'hA01D: data_out = 8'h83;
                    16'hA01E: data_out = 8'h82;
                    16'hA01F: data_out = 8'h81;
                    16'hA020: data_out = 8'h0;
                    16'hA021: data_out = 8'h1;
                    16'hA022: data_out = 8'h2;
                    16'hA023: data_out = 8'h3;
                    16'hA024: data_out = 8'h4;
                    16'hA025: data_out = 8'h5;
                    16'hA026: data_out = 8'h6;
                    16'hA027: data_out = 8'h7;
                    16'hA028: data_out = 8'h8;
                    16'hA029: data_out = 8'h9;
                    16'hA02A: data_out = 8'hA;
                    16'hA02B: data_out = 8'hB;
                    16'hA02C: data_out = 8'hC;
                    16'hA02D: data_out = 8'hD;
                    16'hA02E: data_out = 8'hE;
                    16'hA02F: data_out = 8'hF;
                    16'hA030: data_out = 8'h10;
                    16'hA031: data_out = 8'h11;
                    16'hA032: data_out = 8'h12;
                    16'hA033: data_out = 8'h13;
                    16'hA034: data_out = 8'h14;
                    16'hA035: data_out = 8'h15;
                    16'hA036: data_out = 8'h16;
                    16'hA037: data_out = 8'h17;
                    16'hA038: data_out = 8'h18;
                    16'hA039: data_out = 8'h19;
                    16'hA03A: data_out = 8'h1A;
                    16'hA03B: data_out = 8'h1B;
                    16'hA03C: data_out = 8'h1C;
                    16'hA03D: data_out = 8'h1D;
                    16'hA03E: data_out = 8'h1E;
                    16'hA03F: data_out = 8'h1F;
                    16'hA040: data_out = 8'h20;
                    16'hA041: data_out = 8'h21;
                    16'hA042: data_out = 8'h22;
                    16'hA043: data_out = 8'h23;
                    16'hA044: data_out = 8'h24;
                    16'hA045: data_out = 8'h25;
                    16'hA046: data_out = 8'h26;
                    16'hA047: data_out = 8'h27;
                    16'hA048: data_out = 8'h28;
                    16'hA049: data_out = 8'h29;
                    16'hA04A: data_out = 8'h2A;
                    16'hA04B: data_out = 8'h2B;
                    16'hA04C: data_out = 8'h2C;
                    16'hA04D: data_out = 8'h2D;
                    16'hA04E: data_out = 8'h2E;
                    16'hA04F: data_out = 8'h2F;
                    16'hA050: data_out = 8'h30;
                    16'hA051: data_out = 8'h31;
                    16'hA052: data_out = 8'h32;
                    16'hA053: data_out = 8'h33;
                    16'hA054: data_out = 8'h34;
                    16'hA055: data_out = 8'h35;
                    16'hA056: data_out = 8'h36;
                    16'hA057: data_out = 8'h37;
                    16'hA058: data_out = 8'h38;
                    16'hA059: data_out = 8'h39;
                    16'hA05A: data_out = 8'h3A;
                    16'hA05B: data_out = 8'h3B;
                    16'hA05C: data_out = 8'h3C;
                    16'hA05D: data_out = 8'h3D;
                    16'hA05E: data_out = 8'h3E;
                    16'hA05F: data_out = 8'h3F;
                    16'hA060: data_out = 8'h40;
                    16'hA061: data_out = 8'h41;
                    16'hA062: data_out = 8'h42;
                    16'hA063: data_out = 8'h43;
                    16'hA064: data_out = 8'h44;
                    16'hA065: data_out = 8'h45;
                    16'hA066: data_out = 8'h46;
                    16'hA067: data_out = 8'h47;
                    16'hA068: data_out = 8'h48;
                    16'hA069: data_out = 8'h49;
                    16'hA06A: data_out = 8'h4A;
                    16'hA06B: data_out = 8'h4B;
                    16'hA06C: data_out = 8'h4C;
                    16'hA06D: data_out = 8'h4D;
                    16'hA06E: data_out = 8'h4E;
                    16'hA06F: data_out = 8'h4F;
                    16'hA070: data_out = 8'h50;
                    16'hA071: data_out = 8'h51;
                    16'hA072: data_out = 8'h52;
                    16'hA073: data_out = 8'h53;
                    16'hA074: data_out = 8'h54;
                    16'hA075: data_out = 8'h55;
                    16'hA076: data_out = 8'h56;
                    16'hA077: data_out = 8'h57;
                    16'hA078: data_out = 8'h58;
                    16'hA079: data_out = 8'h59;
                    16'hA07A: data_out = 8'h5A;
                    16'hA07B: data_out = 8'h5B;
                    16'hA07C: data_out = 8'h5C;
                    16'hA07D: data_out = 8'h5D;
                    16'hA07E: data_out = 8'h5E;
                    16'hA07F: data_out = 8'h5F;
                    16'hA080: data_out = 8'hA0;
                    16'hA081: data_out = 8'hA1;
                    16'hA082: data_out = 8'hA2;
                    16'hA083: data_out = 8'hA3;
                    16'hA084: data_out = 8'hA4;
                    16'hA085: data_out = 8'hA5;
                    16'hA086: data_out = 8'hA6;
                    16'hA087: data_out = 8'hA7;
                    16'hA088: data_out = 8'hA8;
                    16'hA089: data_out = 8'hA9;
                    16'hA08A: data_out = 8'hAA;
                    16'hA08B: data_out = 8'hAB;
                    16'hA08C: data_out = 8'hAC;
                    16'hA08D: data_out = 8'hAD;
                    16'hA08E: data_out = 8'hAE;
                    16'hA08F: data_out = 8'hAF;
                    16'hA090: data_out = 8'hB0;
                    16'hA091: data_out = 8'hB1;
                    16'hA092: data_out = 8'hB2;
                    16'hA093: data_out = 8'hB3;
                    16'hA094: data_out = 8'hB4;
                    16'hA095: data_out = 8'hB5;
                    16'hA096: data_out = 8'hB6;
                    16'hA097: data_out = 8'hB7;
                    16'hA098: data_out = 8'hB8;
                    16'hA099: data_out = 8'hB9;
                    16'hA09A: data_out = 8'hBA;
                    16'hA09B: data_out = 8'hBB;
                    16'hA09C: data_out = 8'hBC;
                    16'hA09D: data_out = 8'hBD;
                    16'hA09E: data_out = 8'hBE;
                    16'hA09F: data_out = 8'hBF;
                    16'hA0A0: data_out = 8'hC0;
                    16'hA0A1: data_out = 8'hC1;
                    16'hA0A2: data_out = 8'hC2;
                    16'hA0A3: data_out = 8'hC3;
                    16'hA0A4: data_out = 8'hC4;
                    16'hA0A5: data_out = 8'hC5;
                    16'hA0A6: data_out = 8'hC6;
                    16'hA0A7: data_out = 8'hC7;
                    16'hA0A8: data_out = 8'hC8;
                    16'hA0A9: data_out = 8'hC9;
                    16'hA0AA: data_out = 8'hCA;
                    16'hA0AB: data_out = 8'hCB;
                    16'hA0AC: data_out = 8'hCC;
                    16'hA0AD: data_out = 8'hCD;
                    16'hA0AE: data_out = 8'hCE;
                    16'hA0AF: data_out = 8'hCF;
                    16'hA0B0: data_out = 8'hD0;
                    16'hA0B1: data_out = 8'hD1;
                    16'hA0B2: data_out = 8'hD2;
                    16'hA0B3: data_out = 8'hD3;
                    16'hA0B4: data_out = 8'hD4;
                    16'hA0B5: data_out = 8'hD5;
                    16'hA0B6: data_out = 8'hD6;
                    16'hA0B7: data_out = 8'hD7;
                    16'hA0B8: data_out = 8'hD8;
                    16'hA0B9: data_out = 8'hD9;
                    16'hA0BA: data_out = 8'hDA;
                    16'hA0BB: data_out = 8'hDB;
                    16'hA0BC: data_out = 8'hDC;
                    16'hA0BD: data_out = 8'hDD;
                    16'hA0BE: data_out = 8'hDE;
                    16'hA0BF: data_out = 8'hDF;
                    16'hA0C0: data_out = 8'hE0;
                    16'hA0C1: data_out = 8'hE1;
                    16'hA0C2: data_out = 8'hE2;
                    16'hA0C3: data_out = 8'hE3;
                    16'hA0C4: data_out = 8'hE4;
                    16'hA0C5: data_out = 8'hE5;
                    16'hA0C6: data_out = 8'hE6;
                    16'hA0C7: data_out = 8'hE7;
                    16'hA0C8: data_out = 8'hE8;
                    16'hA0C9: data_out = 8'hE9;
                    16'hA0CA: data_out = 8'hEA;
                    16'hA0CB: data_out = 8'hEB;
                    16'hA0CC: data_out = 8'hEC;
                    16'hA0CD: data_out = 8'hED;
                    16'hA0CE: data_out = 8'hEE;
                    16'hA0CF: data_out = 8'hEF;
                    16'hA0D0: data_out = 8'hF0;
                    16'hA0D1: data_out = 8'hF1;
                    16'hA0D2: data_out = 8'hF2;
                    16'hA0D3: data_out = 8'hF3;
                    16'hA0D4: data_out = 8'hF4;
                    16'hA0D5: data_out = 8'hF5;
                    16'hA0D6: data_out = 8'hF6;
                    16'hA0D7: data_out = 8'hF7;
                    16'hA0D8: data_out = 8'hF8;
                    16'hA0D9: data_out = 8'hF9;
                    16'hA0DA: data_out = 8'hFA;
                    16'hA0DB: data_out = 8'hFB;
                    16'hA0DC: data_out = 8'hFC;
                    16'hA0DD: data_out = 8'hFD;
                    16'hA0DE: data_out = 8'hFE;
                    16'hA0DF: data_out = 8'hFF;
                    16'hA0E0: data_out = 8'h80;
                    16'hA0E1: data_out = 8'h81;
                    16'hA0E2: data_out = 8'h82;
                    16'hA0E3: data_out = 8'h83;
                    16'hA0E4: data_out = 8'h84;
                    16'hA0E5: data_out = 8'h85;
                    16'hA0E6: data_out = 8'h86;
                    16'hA0E7: data_out = 8'h87;
                    16'hA0E8: data_out = 8'h88;
                    16'hA0E9: data_out = 8'h89;
                    16'hA0EA: data_out = 8'h8A;
                    16'hA0EB: data_out = 8'h8B;
                    16'hA0EC: data_out = 8'h8C;
                    16'hA0ED: data_out = 8'h8D;
                    16'hA0EE: data_out = 8'h8E;
                    16'hA0EF: data_out = 8'h8F;
                    16'hA0F0: data_out = 8'h90;
                    16'hA0F1: data_out = 8'h91;
                    16'hA0F2: data_out = 8'h92;
                    16'hA0F3: data_out = 8'h93;
                    16'hA0F4: data_out = 8'h94;
                    16'hA0F5: data_out = 8'h95;
                    16'hA0F6: data_out = 8'h96;
                    16'hA0F7: data_out = 8'h97;
                    16'hA0F8: data_out = 8'h98;
                    16'hA0F9: data_out = 8'h99;
                    16'hA0FA: data_out = 8'h9A;
                    16'hA0FB: data_out = 8'h9B;
                    16'hA0FC: data_out = 8'h9C;
                    16'hA0FD: data_out = 8'h9D;
                    16'hA0FE: data_out = 8'h9E;
                    16'hA0FF: data_out = 8'h9F;
                    16'hA100: data_out = 8'hA1;
                    16'hA101: data_out = 8'hA0;
                    16'hA102: data_out = 8'h9F;
                    16'hA103: data_out = 8'h9E;
                    16'hA104: data_out = 8'h9D;
                    16'hA105: data_out = 8'h9C;
                    16'hA106: data_out = 8'h9B;
                    16'hA107: data_out = 8'h9A;
                    16'hA108: data_out = 8'h99;
                    16'hA109: data_out = 8'h98;
                    16'hA10A: data_out = 8'h97;
                    16'hA10B: data_out = 8'h96;
                    16'hA10C: data_out = 8'h95;
                    16'hA10D: data_out = 8'h94;
                    16'hA10E: data_out = 8'h93;
                    16'hA10F: data_out = 8'h92;
                    16'hA110: data_out = 8'h91;
                    16'hA111: data_out = 8'h90;
                    16'hA112: data_out = 8'h8F;
                    16'hA113: data_out = 8'h8E;
                    16'hA114: data_out = 8'h8D;
                    16'hA115: data_out = 8'h8C;
                    16'hA116: data_out = 8'h8B;
                    16'hA117: data_out = 8'h8A;
                    16'hA118: data_out = 8'h89;
                    16'hA119: data_out = 8'h88;
                    16'hA11A: data_out = 8'h87;
                    16'hA11B: data_out = 8'h86;
                    16'hA11C: data_out = 8'h85;
                    16'hA11D: data_out = 8'h84;
                    16'hA11E: data_out = 8'h83;
                    16'hA11F: data_out = 8'h82;
                    16'hA120: data_out = 8'h81;
                    16'hA121: data_out = 8'h0;
                    16'hA122: data_out = 8'h1;
                    16'hA123: data_out = 8'h2;
                    16'hA124: data_out = 8'h3;
                    16'hA125: data_out = 8'h4;
                    16'hA126: data_out = 8'h5;
                    16'hA127: data_out = 8'h6;
                    16'hA128: data_out = 8'h7;
                    16'hA129: data_out = 8'h8;
                    16'hA12A: data_out = 8'h9;
                    16'hA12B: data_out = 8'hA;
                    16'hA12C: data_out = 8'hB;
                    16'hA12D: data_out = 8'hC;
                    16'hA12E: data_out = 8'hD;
                    16'hA12F: data_out = 8'hE;
                    16'hA130: data_out = 8'hF;
                    16'hA131: data_out = 8'h10;
                    16'hA132: data_out = 8'h11;
                    16'hA133: data_out = 8'h12;
                    16'hA134: data_out = 8'h13;
                    16'hA135: data_out = 8'h14;
                    16'hA136: data_out = 8'h15;
                    16'hA137: data_out = 8'h16;
                    16'hA138: data_out = 8'h17;
                    16'hA139: data_out = 8'h18;
                    16'hA13A: data_out = 8'h19;
                    16'hA13B: data_out = 8'h1A;
                    16'hA13C: data_out = 8'h1B;
                    16'hA13D: data_out = 8'h1C;
                    16'hA13E: data_out = 8'h1D;
                    16'hA13F: data_out = 8'h1E;
                    16'hA140: data_out = 8'h1F;
                    16'hA141: data_out = 8'h20;
                    16'hA142: data_out = 8'h21;
                    16'hA143: data_out = 8'h22;
                    16'hA144: data_out = 8'h23;
                    16'hA145: data_out = 8'h24;
                    16'hA146: data_out = 8'h25;
                    16'hA147: data_out = 8'h26;
                    16'hA148: data_out = 8'h27;
                    16'hA149: data_out = 8'h28;
                    16'hA14A: data_out = 8'h29;
                    16'hA14B: data_out = 8'h2A;
                    16'hA14C: data_out = 8'h2B;
                    16'hA14D: data_out = 8'h2C;
                    16'hA14E: data_out = 8'h2D;
                    16'hA14F: data_out = 8'h2E;
                    16'hA150: data_out = 8'h2F;
                    16'hA151: data_out = 8'h30;
                    16'hA152: data_out = 8'h31;
                    16'hA153: data_out = 8'h32;
                    16'hA154: data_out = 8'h33;
                    16'hA155: data_out = 8'h34;
                    16'hA156: data_out = 8'h35;
                    16'hA157: data_out = 8'h36;
                    16'hA158: data_out = 8'h37;
                    16'hA159: data_out = 8'h38;
                    16'hA15A: data_out = 8'h39;
                    16'hA15B: data_out = 8'h3A;
                    16'hA15C: data_out = 8'h3B;
                    16'hA15D: data_out = 8'h3C;
                    16'hA15E: data_out = 8'h3D;
                    16'hA15F: data_out = 8'h3E;
                    16'hA160: data_out = 8'h3F;
                    16'hA161: data_out = 8'h40;
                    16'hA162: data_out = 8'h41;
                    16'hA163: data_out = 8'h42;
                    16'hA164: data_out = 8'h43;
                    16'hA165: data_out = 8'h44;
                    16'hA166: data_out = 8'h45;
                    16'hA167: data_out = 8'h46;
                    16'hA168: data_out = 8'h47;
                    16'hA169: data_out = 8'h48;
                    16'hA16A: data_out = 8'h49;
                    16'hA16B: data_out = 8'h4A;
                    16'hA16C: data_out = 8'h4B;
                    16'hA16D: data_out = 8'h4C;
                    16'hA16E: data_out = 8'h4D;
                    16'hA16F: data_out = 8'h4E;
                    16'hA170: data_out = 8'h4F;
                    16'hA171: data_out = 8'h50;
                    16'hA172: data_out = 8'h51;
                    16'hA173: data_out = 8'h52;
                    16'hA174: data_out = 8'h53;
                    16'hA175: data_out = 8'h54;
                    16'hA176: data_out = 8'h55;
                    16'hA177: data_out = 8'h56;
                    16'hA178: data_out = 8'h57;
                    16'hA179: data_out = 8'h58;
                    16'hA17A: data_out = 8'h59;
                    16'hA17B: data_out = 8'h5A;
                    16'hA17C: data_out = 8'h5B;
                    16'hA17D: data_out = 8'h5C;
                    16'hA17E: data_out = 8'h5D;
                    16'hA17F: data_out = 8'h5E;
                    16'hA180: data_out = 8'hA1;
                    16'hA181: data_out = 8'hA2;
                    16'hA182: data_out = 8'hA3;
                    16'hA183: data_out = 8'hA4;
                    16'hA184: data_out = 8'hA5;
                    16'hA185: data_out = 8'hA6;
                    16'hA186: data_out = 8'hA7;
                    16'hA187: data_out = 8'hA8;
                    16'hA188: data_out = 8'hA9;
                    16'hA189: data_out = 8'hAA;
                    16'hA18A: data_out = 8'hAB;
                    16'hA18B: data_out = 8'hAC;
                    16'hA18C: data_out = 8'hAD;
                    16'hA18D: data_out = 8'hAE;
                    16'hA18E: data_out = 8'hAF;
                    16'hA18F: data_out = 8'hB0;
                    16'hA190: data_out = 8'hB1;
                    16'hA191: data_out = 8'hB2;
                    16'hA192: data_out = 8'hB3;
                    16'hA193: data_out = 8'hB4;
                    16'hA194: data_out = 8'hB5;
                    16'hA195: data_out = 8'hB6;
                    16'hA196: data_out = 8'hB7;
                    16'hA197: data_out = 8'hB8;
                    16'hA198: data_out = 8'hB9;
                    16'hA199: data_out = 8'hBA;
                    16'hA19A: data_out = 8'hBB;
                    16'hA19B: data_out = 8'hBC;
                    16'hA19C: data_out = 8'hBD;
                    16'hA19D: data_out = 8'hBE;
                    16'hA19E: data_out = 8'hBF;
                    16'hA19F: data_out = 8'hC0;
                    16'hA1A0: data_out = 8'hC1;
                    16'hA1A1: data_out = 8'hC2;
                    16'hA1A2: data_out = 8'hC3;
                    16'hA1A3: data_out = 8'hC4;
                    16'hA1A4: data_out = 8'hC5;
                    16'hA1A5: data_out = 8'hC6;
                    16'hA1A6: data_out = 8'hC7;
                    16'hA1A7: data_out = 8'hC8;
                    16'hA1A8: data_out = 8'hC9;
                    16'hA1A9: data_out = 8'hCA;
                    16'hA1AA: data_out = 8'hCB;
                    16'hA1AB: data_out = 8'hCC;
                    16'hA1AC: data_out = 8'hCD;
                    16'hA1AD: data_out = 8'hCE;
                    16'hA1AE: data_out = 8'hCF;
                    16'hA1AF: data_out = 8'hD0;
                    16'hA1B0: data_out = 8'hD1;
                    16'hA1B1: data_out = 8'hD2;
                    16'hA1B2: data_out = 8'hD3;
                    16'hA1B3: data_out = 8'hD4;
                    16'hA1B4: data_out = 8'hD5;
                    16'hA1B5: data_out = 8'hD6;
                    16'hA1B6: data_out = 8'hD7;
                    16'hA1B7: data_out = 8'hD8;
                    16'hA1B8: data_out = 8'hD9;
                    16'hA1B9: data_out = 8'hDA;
                    16'hA1BA: data_out = 8'hDB;
                    16'hA1BB: data_out = 8'hDC;
                    16'hA1BC: data_out = 8'hDD;
                    16'hA1BD: data_out = 8'hDE;
                    16'hA1BE: data_out = 8'hDF;
                    16'hA1BF: data_out = 8'hE0;
                    16'hA1C0: data_out = 8'hE1;
                    16'hA1C1: data_out = 8'hE2;
                    16'hA1C2: data_out = 8'hE3;
                    16'hA1C3: data_out = 8'hE4;
                    16'hA1C4: data_out = 8'hE5;
                    16'hA1C5: data_out = 8'hE6;
                    16'hA1C6: data_out = 8'hE7;
                    16'hA1C7: data_out = 8'hE8;
                    16'hA1C8: data_out = 8'hE9;
                    16'hA1C9: data_out = 8'hEA;
                    16'hA1CA: data_out = 8'hEB;
                    16'hA1CB: data_out = 8'hEC;
                    16'hA1CC: data_out = 8'hED;
                    16'hA1CD: data_out = 8'hEE;
                    16'hA1CE: data_out = 8'hEF;
                    16'hA1CF: data_out = 8'hF0;
                    16'hA1D0: data_out = 8'hF1;
                    16'hA1D1: data_out = 8'hF2;
                    16'hA1D2: data_out = 8'hF3;
                    16'hA1D3: data_out = 8'hF4;
                    16'hA1D4: data_out = 8'hF5;
                    16'hA1D5: data_out = 8'hF6;
                    16'hA1D6: data_out = 8'hF7;
                    16'hA1D7: data_out = 8'hF8;
                    16'hA1D8: data_out = 8'hF9;
                    16'hA1D9: data_out = 8'hFA;
                    16'hA1DA: data_out = 8'hFB;
                    16'hA1DB: data_out = 8'hFC;
                    16'hA1DC: data_out = 8'hFD;
                    16'hA1DD: data_out = 8'hFE;
                    16'hA1DE: data_out = 8'hFF;
                    16'hA1DF: data_out = 8'h80;
                    16'hA1E0: data_out = 8'h81;
                    16'hA1E1: data_out = 8'h82;
                    16'hA1E2: data_out = 8'h83;
                    16'hA1E3: data_out = 8'h84;
                    16'hA1E4: data_out = 8'h85;
                    16'hA1E5: data_out = 8'h86;
                    16'hA1E6: data_out = 8'h87;
                    16'hA1E7: data_out = 8'h88;
                    16'hA1E8: data_out = 8'h89;
                    16'hA1E9: data_out = 8'h8A;
                    16'hA1EA: data_out = 8'h8B;
                    16'hA1EB: data_out = 8'h8C;
                    16'hA1EC: data_out = 8'h8D;
                    16'hA1ED: data_out = 8'h8E;
                    16'hA1EE: data_out = 8'h8F;
                    16'hA1EF: data_out = 8'h90;
                    16'hA1F0: data_out = 8'h91;
                    16'hA1F1: data_out = 8'h92;
                    16'hA1F2: data_out = 8'h93;
                    16'hA1F3: data_out = 8'h94;
                    16'hA1F4: data_out = 8'h95;
                    16'hA1F5: data_out = 8'h96;
                    16'hA1F6: data_out = 8'h97;
                    16'hA1F7: data_out = 8'h98;
                    16'hA1F8: data_out = 8'h99;
                    16'hA1F9: data_out = 8'h9A;
                    16'hA1FA: data_out = 8'h9B;
                    16'hA1FB: data_out = 8'h9C;
                    16'hA1FC: data_out = 8'h9D;
                    16'hA1FD: data_out = 8'h9E;
                    16'hA1FE: data_out = 8'h9F;
                    16'hA1FF: data_out = 8'hA0;
                    16'hA200: data_out = 8'hA2;
                    16'hA201: data_out = 8'hA1;
                    16'hA202: data_out = 8'hA0;
                    16'hA203: data_out = 8'h9F;
                    16'hA204: data_out = 8'h9E;
                    16'hA205: data_out = 8'h9D;
                    16'hA206: data_out = 8'h9C;
                    16'hA207: data_out = 8'h9B;
                    16'hA208: data_out = 8'h9A;
                    16'hA209: data_out = 8'h99;
                    16'hA20A: data_out = 8'h98;
                    16'hA20B: data_out = 8'h97;
                    16'hA20C: data_out = 8'h96;
                    16'hA20D: data_out = 8'h95;
                    16'hA20E: data_out = 8'h94;
                    16'hA20F: data_out = 8'h93;
                    16'hA210: data_out = 8'h92;
                    16'hA211: data_out = 8'h91;
                    16'hA212: data_out = 8'h90;
                    16'hA213: data_out = 8'h8F;
                    16'hA214: data_out = 8'h8E;
                    16'hA215: data_out = 8'h8D;
                    16'hA216: data_out = 8'h8C;
                    16'hA217: data_out = 8'h8B;
                    16'hA218: data_out = 8'h8A;
                    16'hA219: data_out = 8'h89;
                    16'hA21A: data_out = 8'h88;
                    16'hA21B: data_out = 8'h87;
                    16'hA21C: data_out = 8'h86;
                    16'hA21D: data_out = 8'h85;
                    16'hA21E: data_out = 8'h84;
                    16'hA21F: data_out = 8'h83;
                    16'hA220: data_out = 8'h82;
                    16'hA221: data_out = 8'h81;
                    16'hA222: data_out = 8'h0;
                    16'hA223: data_out = 8'h1;
                    16'hA224: data_out = 8'h2;
                    16'hA225: data_out = 8'h3;
                    16'hA226: data_out = 8'h4;
                    16'hA227: data_out = 8'h5;
                    16'hA228: data_out = 8'h6;
                    16'hA229: data_out = 8'h7;
                    16'hA22A: data_out = 8'h8;
                    16'hA22B: data_out = 8'h9;
                    16'hA22C: data_out = 8'hA;
                    16'hA22D: data_out = 8'hB;
                    16'hA22E: data_out = 8'hC;
                    16'hA22F: data_out = 8'hD;
                    16'hA230: data_out = 8'hE;
                    16'hA231: data_out = 8'hF;
                    16'hA232: data_out = 8'h10;
                    16'hA233: data_out = 8'h11;
                    16'hA234: data_out = 8'h12;
                    16'hA235: data_out = 8'h13;
                    16'hA236: data_out = 8'h14;
                    16'hA237: data_out = 8'h15;
                    16'hA238: data_out = 8'h16;
                    16'hA239: data_out = 8'h17;
                    16'hA23A: data_out = 8'h18;
                    16'hA23B: data_out = 8'h19;
                    16'hA23C: data_out = 8'h1A;
                    16'hA23D: data_out = 8'h1B;
                    16'hA23E: data_out = 8'h1C;
                    16'hA23F: data_out = 8'h1D;
                    16'hA240: data_out = 8'h1E;
                    16'hA241: data_out = 8'h1F;
                    16'hA242: data_out = 8'h20;
                    16'hA243: data_out = 8'h21;
                    16'hA244: data_out = 8'h22;
                    16'hA245: data_out = 8'h23;
                    16'hA246: data_out = 8'h24;
                    16'hA247: data_out = 8'h25;
                    16'hA248: data_out = 8'h26;
                    16'hA249: data_out = 8'h27;
                    16'hA24A: data_out = 8'h28;
                    16'hA24B: data_out = 8'h29;
                    16'hA24C: data_out = 8'h2A;
                    16'hA24D: data_out = 8'h2B;
                    16'hA24E: data_out = 8'h2C;
                    16'hA24F: data_out = 8'h2D;
                    16'hA250: data_out = 8'h2E;
                    16'hA251: data_out = 8'h2F;
                    16'hA252: data_out = 8'h30;
                    16'hA253: data_out = 8'h31;
                    16'hA254: data_out = 8'h32;
                    16'hA255: data_out = 8'h33;
                    16'hA256: data_out = 8'h34;
                    16'hA257: data_out = 8'h35;
                    16'hA258: data_out = 8'h36;
                    16'hA259: data_out = 8'h37;
                    16'hA25A: data_out = 8'h38;
                    16'hA25B: data_out = 8'h39;
                    16'hA25C: data_out = 8'h3A;
                    16'hA25D: data_out = 8'h3B;
                    16'hA25E: data_out = 8'h3C;
                    16'hA25F: data_out = 8'h3D;
                    16'hA260: data_out = 8'h3E;
                    16'hA261: data_out = 8'h3F;
                    16'hA262: data_out = 8'h40;
                    16'hA263: data_out = 8'h41;
                    16'hA264: data_out = 8'h42;
                    16'hA265: data_out = 8'h43;
                    16'hA266: data_out = 8'h44;
                    16'hA267: data_out = 8'h45;
                    16'hA268: data_out = 8'h46;
                    16'hA269: data_out = 8'h47;
                    16'hA26A: data_out = 8'h48;
                    16'hA26B: data_out = 8'h49;
                    16'hA26C: data_out = 8'h4A;
                    16'hA26D: data_out = 8'h4B;
                    16'hA26E: data_out = 8'h4C;
                    16'hA26F: data_out = 8'h4D;
                    16'hA270: data_out = 8'h4E;
                    16'hA271: data_out = 8'h4F;
                    16'hA272: data_out = 8'h50;
                    16'hA273: data_out = 8'h51;
                    16'hA274: data_out = 8'h52;
                    16'hA275: data_out = 8'h53;
                    16'hA276: data_out = 8'h54;
                    16'hA277: data_out = 8'h55;
                    16'hA278: data_out = 8'h56;
                    16'hA279: data_out = 8'h57;
                    16'hA27A: data_out = 8'h58;
                    16'hA27B: data_out = 8'h59;
                    16'hA27C: data_out = 8'h5A;
                    16'hA27D: data_out = 8'h5B;
                    16'hA27E: data_out = 8'h5C;
                    16'hA27F: data_out = 8'h5D;
                    16'hA280: data_out = 8'hA2;
                    16'hA281: data_out = 8'hA3;
                    16'hA282: data_out = 8'hA4;
                    16'hA283: data_out = 8'hA5;
                    16'hA284: data_out = 8'hA6;
                    16'hA285: data_out = 8'hA7;
                    16'hA286: data_out = 8'hA8;
                    16'hA287: data_out = 8'hA9;
                    16'hA288: data_out = 8'hAA;
                    16'hA289: data_out = 8'hAB;
                    16'hA28A: data_out = 8'hAC;
                    16'hA28B: data_out = 8'hAD;
                    16'hA28C: data_out = 8'hAE;
                    16'hA28D: data_out = 8'hAF;
                    16'hA28E: data_out = 8'hB0;
                    16'hA28F: data_out = 8'hB1;
                    16'hA290: data_out = 8'hB2;
                    16'hA291: data_out = 8'hB3;
                    16'hA292: data_out = 8'hB4;
                    16'hA293: data_out = 8'hB5;
                    16'hA294: data_out = 8'hB6;
                    16'hA295: data_out = 8'hB7;
                    16'hA296: data_out = 8'hB8;
                    16'hA297: data_out = 8'hB9;
                    16'hA298: data_out = 8'hBA;
                    16'hA299: data_out = 8'hBB;
                    16'hA29A: data_out = 8'hBC;
                    16'hA29B: data_out = 8'hBD;
                    16'hA29C: data_out = 8'hBE;
                    16'hA29D: data_out = 8'hBF;
                    16'hA29E: data_out = 8'hC0;
                    16'hA29F: data_out = 8'hC1;
                    16'hA2A0: data_out = 8'hC2;
                    16'hA2A1: data_out = 8'hC3;
                    16'hA2A2: data_out = 8'hC4;
                    16'hA2A3: data_out = 8'hC5;
                    16'hA2A4: data_out = 8'hC6;
                    16'hA2A5: data_out = 8'hC7;
                    16'hA2A6: data_out = 8'hC8;
                    16'hA2A7: data_out = 8'hC9;
                    16'hA2A8: data_out = 8'hCA;
                    16'hA2A9: data_out = 8'hCB;
                    16'hA2AA: data_out = 8'hCC;
                    16'hA2AB: data_out = 8'hCD;
                    16'hA2AC: data_out = 8'hCE;
                    16'hA2AD: data_out = 8'hCF;
                    16'hA2AE: data_out = 8'hD0;
                    16'hA2AF: data_out = 8'hD1;
                    16'hA2B0: data_out = 8'hD2;
                    16'hA2B1: data_out = 8'hD3;
                    16'hA2B2: data_out = 8'hD4;
                    16'hA2B3: data_out = 8'hD5;
                    16'hA2B4: data_out = 8'hD6;
                    16'hA2B5: data_out = 8'hD7;
                    16'hA2B6: data_out = 8'hD8;
                    16'hA2B7: data_out = 8'hD9;
                    16'hA2B8: data_out = 8'hDA;
                    16'hA2B9: data_out = 8'hDB;
                    16'hA2BA: data_out = 8'hDC;
                    16'hA2BB: data_out = 8'hDD;
                    16'hA2BC: data_out = 8'hDE;
                    16'hA2BD: data_out = 8'hDF;
                    16'hA2BE: data_out = 8'hE0;
                    16'hA2BF: data_out = 8'hE1;
                    16'hA2C0: data_out = 8'hE2;
                    16'hA2C1: data_out = 8'hE3;
                    16'hA2C2: data_out = 8'hE4;
                    16'hA2C3: data_out = 8'hE5;
                    16'hA2C4: data_out = 8'hE6;
                    16'hA2C5: data_out = 8'hE7;
                    16'hA2C6: data_out = 8'hE8;
                    16'hA2C7: data_out = 8'hE9;
                    16'hA2C8: data_out = 8'hEA;
                    16'hA2C9: data_out = 8'hEB;
                    16'hA2CA: data_out = 8'hEC;
                    16'hA2CB: data_out = 8'hED;
                    16'hA2CC: data_out = 8'hEE;
                    16'hA2CD: data_out = 8'hEF;
                    16'hA2CE: data_out = 8'hF0;
                    16'hA2CF: data_out = 8'hF1;
                    16'hA2D0: data_out = 8'hF2;
                    16'hA2D1: data_out = 8'hF3;
                    16'hA2D2: data_out = 8'hF4;
                    16'hA2D3: data_out = 8'hF5;
                    16'hA2D4: data_out = 8'hF6;
                    16'hA2D5: data_out = 8'hF7;
                    16'hA2D6: data_out = 8'hF8;
                    16'hA2D7: data_out = 8'hF9;
                    16'hA2D8: data_out = 8'hFA;
                    16'hA2D9: data_out = 8'hFB;
                    16'hA2DA: data_out = 8'hFC;
                    16'hA2DB: data_out = 8'hFD;
                    16'hA2DC: data_out = 8'hFE;
                    16'hA2DD: data_out = 8'hFF;
                    16'hA2DE: data_out = 8'h80;
                    16'hA2DF: data_out = 8'h81;
                    16'hA2E0: data_out = 8'h82;
                    16'hA2E1: data_out = 8'h83;
                    16'hA2E2: data_out = 8'h84;
                    16'hA2E3: data_out = 8'h85;
                    16'hA2E4: data_out = 8'h86;
                    16'hA2E5: data_out = 8'h87;
                    16'hA2E6: data_out = 8'h88;
                    16'hA2E7: data_out = 8'h89;
                    16'hA2E8: data_out = 8'h8A;
                    16'hA2E9: data_out = 8'h8B;
                    16'hA2EA: data_out = 8'h8C;
                    16'hA2EB: data_out = 8'h8D;
                    16'hA2EC: data_out = 8'h8E;
                    16'hA2ED: data_out = 8'h8F;
                    16'hA2EE: data_out = 8'h90;
                    16'hA2EF: data_out = 8'h91;
                    16'hA2F0: data_out = 8'h92;
                    16'hA2F1: data_out = 8'h93;
                    16'hA2F2: data_out = 8'h94;
                    16'hA2F3: data_out = 8'h95;
                    16'hA2F4: data_out = 8'h96;
                    16'hA2F5: data_out = 8'h97;
                    16'hA2F6: data_out = 8'h98;
                    16'hA2F7: data_out = 8'h99;
                    16'hA2F8: data_out = 8'h9A;
                    16'hA2F9: data_out = 8'h9B;
                    16'hA2FA: data_out = 8'h9C;
                    16'hA2FB: data_out = 8'h9D;
                    16'hA2FC: data_out = 8'h9E;
                    16'hA2FD: data_out = 8'h9F;
                    16'hA2FE: data_out = 8'hA0;
                    16'hA2FF: data_out = 8'hA1;
                    16'hA300: data_out = 8'hA3;
                    16'hA301: data_out = 8'hA2;
                    16'hA302: data_out = 8'hA1;
                    16'hA303: data_out = 8'hA0;
                    16'hA304: data_out = 8'h9F;
                    16'hA305: data_out = 8'h9E;
                    16'hA306: data_out = 8'h9D;
                    16'hA307: data_out = 8'h9C;
                    16'hA308: data_out = 8'h9B;
                    16'hA309: data_out = 8'h9A;
                    16'hA30A: data_out = 8'h99;
                    16'hA30B: data_out = 8'h98;
                    16'hA30C: data_out = 8'h97;
                    16'hA30D: data_out = 8'h96;
                    16'hA30E: data_out = 8'h95;
                    16'hA30F: data_out = 8'h94;
                    16'hA310: data_out = 8'h93;
                    16'hA311: data_out = 8'h92;
                    16'hA312: data_out = 8'h91;
                    16'hA313: data_out = 8'h90;
                    16'hA314: data_out = 8'h8F;
                    16'hA315: data_out = 8'h8E;
                    16'hA316: data_out = 8'h8D;
                    16'hA317: data_out = 8'h8C;
                    16'hA318: data_out = 8'h8B;
                    16'hA319: data_out = 8'h8A;
                    16'hA31A: data_out = 8'h89;
                    16'hA31B: data_out = 8'h88;
                    16'hA31C: data_out = 8'h87;
                    16'hA31D: data_out = 8'h86;
                    16'hA31E: data_out = 8'h85;
                    16'hA31F: data_out = 8'h84;
                    16'hA320: data_out = 8'h83;
                    16'hA321: data_out = 8'h82;
                    16'hA322: data_out = 8'h81;
                    16'hA323: data_out = 8'h0;
                    16'hA324: data_out = 8'h1;
                    16'hA325: data_out = 8'h2;
                    16'hA326: data_out = 8'h3;
                    16'hA327: data_out = 8'h4;
                    16'hA328: data_out = 8'h5;
                    16'hA329: data_out = 8'h6;
                    16'hA32A: data_out = 8'h7;
                    16'hA32B: data_out = 8'h8;
                    16'hA32C: data_out = 8'h9;
                    16'hA32D: data_out = 8'hA;
                    16'hA32E: data_out = 8'hB;
                    16'hA32F: data_out = 8'hC;
                    16'hA330: data_out = 8'hD;
                    16'hA331: data_out = 8'hE;
                    16'hA332: data_out = 8'hF;
                    16'hA333: data_out = 8'h10;
                    16'hA334: data_out = 8'h11;
                    16'hA335: data_out = 8'h12;
                    16'hA336: data_out = 8'h13;
                    16'hA337: data_out = 8'h14;
                    16'hA338: data_out = 8'h15;
                    16'hA339: data_out = 8'h16;
                    16'hA33A: data_out = 8'h17;
                    16'hA33B: data_out = 8'h18;
                    16'hA33C: data_out = 8'h19;
                    16'hA33D: data_out = 8'h1A;
                    16'hA33E: data_out = 8'h1B;
                    16'hA33F: data_out = 8'h1C;
                    16'hA340: data_out = 8'h1D;
                    16'hA341: data_out = 8'h1E;
                    16'hA342: data_out = 8'h1F;
                    16'hA343: data_out = 8'h20;
                    16'hA344: data_out = 8'h21;
                    16'hA345: data_out = 8'h22;
                    16'hA346: data_out = 8'h23;
                    16'hA347: data_out = 8'h24;
                    16'hA348: data_out = 8'h25;
                    16'hA349: data_out = 8'h26;
                    16'hA34A: data_out = 8'h27;
                    16'hA34B: data_out = 8'h28;
                    16'hA34C: data_out = 8'h29;
                    16'hA34D: data_out = 8'h2A;
                    16'hA34E: data_out = 8'h2B;
                    16'hA34F: data_out = 8'h2C;
                    16'hA350: data_out = 8'h2D;
                    16'hA351: data_out = 8'h2E;
                    16'hA352: data_out = 8'h2F;
                    16'hA353: data_out = 8'h30;
                    16'hA354: data_out = 8'h31;
                    16'hA355: data_out = 8'h32;
                    16'hA356: data_out = 8'h33;
                    16'hA357: data_out = 8'h34;
                    16'hA358: data_out = 8'h35;
                    16'hA359: data_out = 8'h36;
                    16'hA35A: data_out = 8'h37;
                    16'hA35B: data_out = 8'h38;
                    16'hA35C: data_out = 8'h39;
                    16'hA35D: data_out = 8'h3A;
                    16'hA35E: data_out = 8'h3B;
                    16'hA35F: data_out = 8'h3C;
                    16'hA360: data_out = 8'h3D;
                    16'hA361: data_out = 8'h3E;
                    16'hA362: data_out = 8'h3F;
                    16'hA363: data_out = 8'h40;
                    16'hA364: data_out = 8'h41;
                    16'hA365: data_out = 8'h42;
                    16'hA366: data_out = 8'h43;
                    16'hA367: data_out = 8'h44;
                    16'hA368: data_out = 8'h45;
                    16'hA369: data_out = 8'h46;
                    16'hA36A: data_out = 8'h47;
                    16'hA36B: data_out = 8'h48;
                    16'hA36C: data_out = 8'h49;
                    16'hA36D: data_out = 8'h4A;
                    16'hA36E: data_out = 8'h4B;
                    16'hA36F: data_out = 8'h4C;
                    16'hA370: data_out = 8'h4D;
                    16'hA371: data_out = 8'h4E;
                    16'hA372: data_out = 8'h4F;
                    16'hA373: data_out = 8'h50;
                    16'hA374: data_out = 8'h51;
                    16'hA375: data_out = 8'h52;
                    16'hA376: data_out = 8'h53;
                    16'hA377: data_out = 8'h54;
                    16'hA378: data_out = 8'h55;
                    16'hA379: data_out = 8'h56;
                    16'hA37A: data_out = 8'h57;
                    16'hA37B: data_out = 8'h58;
                    16'hA37C: data_out = 8'h59;
                    16'hA37D: data_out = 8'h5A;
                    16'hA37E: data_out = 8'h5B;
                    16'hA37F: data_out = 8'h5C;
                    16'hA380: data_out = 8'hA3;
                    16'hA381: data_out = 8'hA4;
                    16'hA382: data_out = 8'hA5;
                    16'hA383: data_out = 8'hA6;
                    16'hA384: data_out = 8'hA7;
                    16'hA385: data_out = 8'hA8;
                    16'hA386: data_out = 8'hA9;
                    16'hA387: data_out = 8'hAA;
                    16'hA388: data_out = 8'hAB;
                    16'hA389: data_out = 8'hAC;
                    16'hA38A: data_out = 8'hAD;
                    16'hA38B: data_out = 8'hAE;
                    16'hA38C: data_out = 8'hAF;
                    16'hA38D: data_out = 8'hB0;
                    16'hA38E: data_out = 8'hB1;
                    16'hA38F: data_out = 8'hB2;
                    16'hA390: data_out = 8'hB3;
                    16'hA391: data_out = 8'hB4;
                    16'hA392: data_out = 8'hB5;
                    16'hA393: data_out = 8'hB6;
                    16'hA394: data_out = 8'hB7;
                    16'hA395: data_out = 8'hB8;
                    16'hA396: data_out = 8'hB9;
                    16'hA397: data_out = 8'hBA;
                    16'hA398: data_out = 8'hBB;
                    16'hA399: data_out = 8'hBC;
                    16'hA39A: data_out = 8'hBD;
                    16'hA39B: data_out = 8'hBE;
                    16'hA39C: data_out = 8'hBF;
                    16'hA39D: data_out = 8'hC0;
                    16'hA39E: data_out = 8'hC1;
                    16'hA39F: data_out = 8'hC2;
                    16'hA3A0: data_out = 8'hC3;
                    16'hA3A1: data_out = 8'hC4;
                    16'hA3A2: data_out = 8'hC5;
                    16'hA3A3: data_out = 8'hC6;
                    16'hA3A4: data_out = 8'hC7;
                    16'hA3A5: data_out = 8'hC8;
                    16'hA3A6: data_out = 8'hC9;
                    16'hA3A7: data_out = 8'hCA;
                    16'hA3A8: data_out = 8'hCB;
                    16'hA3A9: data_out = 8'hCC;
                    16'hA3AA: data_out = 8'hCD;
                    16'hA3AB: data_out = 8'hCE;
                    16'hA3AC: data_out = 8'hCF;
                    16'hA3AD: data_out = 8'hD0;
                    16'hA3AE: data_out = 8'hD1;
                    16'hA3AF: data_out = 8'hD2;
                    16'hA3B0: data_out = 8'hD3;
                    16'hA3B1: data_out = 8'hD4;
                    16'hA3B2: data_out = 8'hD5;
                    16'hA3B3: data_out = 8'hD6;
                    16'hA3B4: data_out = 8'hD7;
                    16'hA3B5: data_out = 8'hD8;
                    16'hA3B6: data_out = 8'hD9;
                    16'hA3B7: data_out = 8'hDA;
                    16'hA3B8: data_out = 8'hDB;
                    16'hA3B9: data_out = 8'hDC;
                    16'hA3BA: data_out = 8'hDD;
                    16'hA3BB: data_out = 8'hDE;
                    16'hA3BC: data_out = 8'hDF;
                    16'hA3BD: data_out = 8'hE0;
                    16'hA3BE: data_out = 8'hE1;
                    16'hA3BF: data_out = 8'hE2;
                    16'hA3C0: data_out = 8'hE3;
                    16'hA3C1: data_out = 8'hE4;
                    16'hA3C2: data_out = 8'hE5;
                    16'hA3C3: data_out = 8'hE6;
                    16'hA3C4: data_out = 8'hE7;
                    16'hA3C5: data_out = 8'hE8;
                    16'hA3C6: data_out = 8'hE9;
                    16'hA3C7: data_out = 8'hEA;
                    16'hA3C8: data_out = 8'hEB;
                    16'hA3C9: data_out = 8'hEC;
                    16'hA3CA: data_out = 8'hED;
                    16'hA3CB: data_out = 8'hEE;
                    16'hA3CC: data_out = 8'hEF;
                    16'hA3CD: data_out = 8'hF0;
                    16'hA3CE: data_out = 8'hF1;
                    16'hA3CF: data_out = 8'hF2;
                    16'hA3D0: data_out = 8'hF3;
                    16'hA3D1: data_out = 8'hF4;
                    16'hA3D2: data_out = 8'hF5;
                    16'hA3D3: data_out = 8'hF6;
                    16'hA3D4: data_out = 8'hF7;
                    16'hA3D5: data_out = 8'hF8;
                    16'hA3D6: data_out = 8'hF9;
                    16'hA3D7: data_out = 8'hFA;
                    16'hA3D8: data_out = 8'hFB;
                    16'hA3D9: data_out = 8'hFC;
                    16'hA3DA: data_out = 8'hFD;
                    16'hA3DB: data_out = 8'hFE;
                    16'hA3DC: data_out = 8'hFF;
                    16'hA3DD: data_out = 8'h80;
                    16'hA3DE: data_out = 8'h81;
                    16'hA3DF: data_out = 8'h82;
                    16'hA3E0: data_out = 8'h83;
                    16'hA3E1: data_out = 8'h84;
                    16'hA3E2: data_out = 8'h85;
                    16'hA3E3: data_out = 8'h86;
                    16'hA3E4: data_out = 8'h87;
                    16'hA3E5: data_out = 8'h88;
                    16'hA3E6: data_out = 8'h89;
                    16'hA3E7: data_out = 8'h8A;
                    16'hA3E8: data_out = 8'h8B;
                    16'hA3E9: data_out = 8'h8C;
                    16'hA3EA: data_out = 8'h8D;
                    16'hA3EB: data_out = 8'h8E;
                    16'hA3EC: data_out = 8'h8F;
                    16'hA3ED: data_out = 8'h90;
                    16'hA3EE: data_out = 8'h91;
                    16'hA3EF: data_out = 8'h92;
                    16'hA3F0: data_out = 8'h93;
                    16'hA3F1: data_out = 8'h94;
                    16'hA3F2: data_out = 8'h95;
                    16'hA3F3: data_out = 8'h96;
                    16'hA3F4: data_out = 8'h97;
                    16'hA3F5: data_out = 8'h98;
                    16'hA3F6: data_out = 8'h99;
                    16'hA3F7: data_out = 8'h9A;
                    16'hA3F8: data_out = 8'h9B;
                    16'hA3F9: data_out = 8'h9C;
                    16'hA3FA: data_out = 8'h9D;
                    16'hA3FB: data_out = 8'h9E;
                    16'hA3FC: data_out = 8'h9F;
                    16'hA3FD: data_out = 8'hA0;
                    16'hA3FE: data_out = 8'hA1;
                    16'hA3FF: data_out = 8'hA2;
                    16'hA400: data_out = 8'hA4;
                    16'hA401: data_out = 8'hA3;
                    16'hA402: data_out = 8'hA2;
                    16'hA403: data_out = 8'hA1;
                    16'hA404: data_out = 8'hA0;
                    16'hA405: data_out = 8'h9F;
                    16'hA406: data_out = 8'h9E;
                    16'hA407: data_out = 8'h9D;
                    16'hA408: data_out = 8'h9C;
                    16'hA409: data_out = 8'h9B;
                    16'hA40A: data_out = 8'h9A;
                    16'hA40B: data_out = 8'h99;
                    16'hA40C: data_out = 8'h98;
                    16'hA40D: data_out = 8'h97;
                    16'hA40E: data_out = 8'h96;
                    16'hA40F: data_out = 8'h95;
                    16'hA410: data_out = 8'h94;
                    16'hA411: data_out = 8'h93;
                    16'hA412: data_out = 8'h92;
                    16'hA413: data_out = 8'h91;
                    16'hA414: data_out = 8'h90;
                    16'hA415: data_out = 8'h8F;
                    16'hA416: data_out = 8'h8E;
                    16'hA417: data_out = 8'h8D;
                    16'hA418: data_out = 8'h8C;
                    16'hA419: data_out = 8'h8B;
                    16'hA41A: data_out = 8'h8A;
                    16'hA41B: data_out = 8'h89;
                    16'hA41C: data_out = 8'h88;
                    16'hA41D: data_out = 8'h87;
                    16'hA41E: data_out = 8'h86;
                    16'hA41F: data_out = 8'h85;
                    16'hA420: data_out = 8'h84;
                    16'hA421: data_out = 8'h83;
                    16'hA422: data_out = 8'h82;
                    16'hA423: data_out = 8'h81;
                    16'hA424: data_out = 8'h0;
                    16'hA425: data_out = 8'h1;
                    16'hA426: data_out = 8'h2;
                    16'hA427: data_out = 8'h3;
                    16'hA428: data_out = 8'h4;
                    16'hA429: data_out = 8'h5;
                    16'hA42A: data_out = 8'h6;
                    16'hA42B: data_out = 8'h7;
                    16'hA42C: data_out = 8'h8;
                    16'hA42D: data_out = 8'h9;
                    16'hA42E: data_out = 8'hA;
                    16'hA42F: data_out = 8'hB;
                    16'hA430: data_out = 8'hC;
                    16'hA431: data_out = 8'hD;
                    16'hA432: data_out = 8'hE;
                    16'hA433: data_out = 8'hF;
                    16'hA434: data_out = 8'h10;
                    16'hA435: data_out = 8'h11;
                    16'hA436: data_out = 8'h12;
                    16'hA437: data_out = 8'h13;
                    16'hA438: data_out = 8'h14;
                    16'hA439: data_out = 8'h15;
                    16'hA43A: data_out = 8'h16;
                    16'hA43B: data_out = 8'h17;
                    16'hA43C: data_out = 8'h18;
                    16'hA43D: data_out = 8'h19;
                    16'hA43E: data_out = 8'h1A;
                    16'hA43F: data_out = 8'h1B;
                    16'hA440: data_out = 8'h1C;
                    16'hA441: data_out = 8'h1D;
                    16'hA442: data_out = 8'h1E;
                    16'hA443: data_out = 8'h1F;
                    16'hA444: data_out = 8'h20;
                    16'hA445: data_out = 8'h21;
                    16'hA446: data_out = 8'h22;
                    16'hA447: data_out = 8'h23;
                    16'hA448: data_out = 8'h24;
                    16'hA449: data_out = 8'h25;
                    16'hA44A: data_out = 8'h26;
                    16'hA44B: data_out = 8'h27;
                    16'hA44C: data_out = 8'h28;
                    16'hA44D: data_out = 8'h29;
                    16'hA44E: data_out = 8'h2A;
                    16'hA44F: data_out = 8'h2B;
                    16'hA450: data_out = 8'h2C;
                    16'hA451: data_out = 8'h2D;
                    16'hA452: data_out = 8'h2E;
                    16'hA453: data_out = 8'h2F;
                    16'hA454: data_out = 8'h30;
                    16'hA455: data_out = 8'h31;
                    16'hA456: data_out = 8'h32;
                    16'hA457: data_out = 8'h33;
                    16'hA458: data_out = 8'h34;
                    16'hA459: data_out = 8'h35;
                    16'hA45A: data_out = 8'h36;
                    16'hA45B: data_out = 8'h37;
                    16'hA45C: data_out = 8'h38;
                    16'hA45D: data_out = 8'h39;
                    16'hA45E: data_out = 8'h3A;
                    16'hA45F: data_out = 8'h3B;
                    16'hA460: data_out = 8'h3C;
                    16'hA461: data_out = 8'h3D;
                    16'hA462: data_out = 8'h3E;
                    16'hA463: data_out = 8'h3F;
                    16'hA464: data_out = 8'h40;
                    16'hA465: data_out = 8'h41;
                    16'hA466: data_out = 8'h42;
                    16'hA467: data_out = 8'h43;
                    16'hA468: data_out = 8'h44;
                    16'hA469: data_out = 8'h45;
                    16'hA46A: data_out = 8'h46;
                    16'hA46B: data_out = 8'h47;
                    16'hA46C: data_out = 8'h48;
                    16'hA46D: data_out = 8'h49;
                    16'hA46E: data_out = 8'h4A;
                    16'hA46F: data_out = 8'h4B;
                    16'hA470: data_out = 8'h4C;
                    16'hA471: data_out = 8'h4D;
                    16'hA472: data_out = 8'h4E;
                    16'hA473: data_out = 8'h4F;
                    16'hA474: data_out = 8'h50;
                    16'hA475: data_out = 8'h51;
                    16'hA476: data_out = 8'h52;
                    16'hA477: data_out = 8'h53;
                    16'hA478: data_out = 8'h54;
                    16'hA479: data_out = 8'h55;
                    16'hA47A: data_out = 8'h56;
                    16'hA47B: data_out = 8'h57;
                    16'hA47C: data_out = 8'h58;
                    16'hA47D: data_out = 8'h59;
                    16'hA47E: data_out = 8'h5A;
                    16'hA47F: data_out = 8'h5B;
                    16'hA480: data_out = 8'hA4;
                    16'hA481: data_out = 8'hA5;
                    16'hA482: data_out = 8'hA6;
                    16'hA483: data_out = 8'hA7;
                    16'hA484: data_out = 8'hA8;
                    16'hA485: data_out = 8'hA9;
                    16'hA486: data_out = 8'hAA;
                    16'hA487: data_out = 8'hAB;
                    16'hA488: data_out = 8'hAC;
                    16'hA489: data_out = 8'hAD;
                    16'hA48A: data_out = 8'hAE;
                    16'hA48B: data_out = 8'hAF;
                    16'hA48C: data_out = 8'hB0;
                    16'hA48D: data_out = 8'hB1;
                    16'hA48E: data_out = 8'hB2;
                    16'hA48F: data_out = 8'hB3;
                    16'hA490: data_out = 8'hB4;
                    16'hA491: data_out = 8'hB5;
                    16'hA492: data_out = 8'hB6;
                    16'hA493: data_out = 8'hB7;
                    16'hA494: data_out = 8'hB8;
                    16'hA495: data_out = 8'hB9;
                    16'hA496: data_out = 8'hBA;
                    16'hA497: data_out = 8'hBB;
                    16'hA498: data_out = 8'hBC;
                    16'hA499: data_out = 8'hBD;
                    16'hA49A: data_out = 8'hBE;
                    16'hA49B: data_out = 8'hBF;
                    16'hA49C: data_out = 8'hC0;
                    16'hA49D: data_out = 8'hC1;
                    16'hA49E: data_out = 8'hC2;
                    16'hA49F: data_out = 8'hC3;
                    16'hA4A0: data_out = 8'hC4;
                    16'hA4A1: data_out = 8'hC5;
                    16'hA4A2: data_out = 8'hC6;
                    16'hA4A3: data_out = 8'hC7;
                    16'hA4A4: data_out = 8'hC8;
                    16'hA4A5: data_out = 8'hC9;
                    16'hA4A6: data_out = 8'hCA;
                    16'hA4A7: data_out = 8'hCB;
                    16'hA4A8: data_out = 8'hCC;
                    16'hA4A9: data_out = 8'hCD;
                    16'hA4AA: data_out = 8'hCE;
                    16'hA4AB: data_out = 8'hCF;
                    16'hA4AC: data_out = 8'hD0;
                    16'hA4AD: data_out = 8'hD1;
                    16'hA4AE: data_out = 8'hD2;
                    16'hA4AF: data_out = 8'hD3;
                    16'hA4B0: data_out = 8'hD4;
                    16'hA4B1: data_out = 8'hD5;
                    16'hA4B2: data_out = 8'hD6;
                    16'hA4B3: data_out = 8'hD7;
                    16'hA4B4: data_out = 8'hD8;
                    16'hA4B5: data_out = 8'hD9;
                    16'hA4B6: data_out = 8'hDA;
                    16'hA4B7: data_out = 8'hDB;
                    16'hA4B8: data_out = 8'hDC;
                    16'hA4B9: data_out = 8'hDD;
                    16'hA4BA: data_out = 8'hDE;
                    16'hA4BB: data_out = 8'hDF;
                    16'hA4BC: data_out = 8'hE0;
                    16'hA4BD: data_out = 8'hE1;
                    16'hA4BE: data_out = 8'hE2;
                    16'hA4BF: data_out = 8'hE3;
                    16'hA4C0: data_out = 8'hE4;
                    16'hA4C1: data_out = 8'hE5;
                    16'hA4C2: data_out = 8'hE6;
                    16'hA4C3: data_out = 8'hE7;
                    16'hA4C4: data_out = 8'hE8;
                    16'hA4C5: data_out = 8'hE9;
                    16'hA4C6: data_out = 8'hEA;
                    16'hA4C7: data_out = 8'hEB;
                    16'hA4C8: data_out = 8'hEC;
                    16'hA4C9: data_out = 8'hED;
                    16'hA4CA: data_out = 8'hEE;
                    16'hA4CB: data_out = 8'hEF;
                    16'hA4CC: data_out = 8'hF0;
                    16'hA4CD: data_out = 8'hF1;
                    16'hA4CE: data_out = 8'hF2;
                    16'hA4CF: data_out = 8'hF3;
                    16'hA4D0: data_out = 8'hF4;
                    16'hA4D1: data_out = 8'hF5;
                    16'hA4D2: data_out = 8'hF6;
                    16'hA4D3: data_out = 8'hF7;
                    16'hA4D4: data_out = 8'hF8;
                    16'hA4D5: data_out = 8'hF9;
                    16'hA4D6: data_out = 8'hFA;
                    16'hA4D7: data_out = 8'hFB;
                    16'hA4D8: data_out = 8'hFC;
                    16'hA4D9: data_out = 8'hFD;
                    16'hA4DA: data_out = 8'hFE;
                    16'hA4DB: data_out = 8'hFF;
                    16'hA4DC: data_out = 8'h80;
                    16'hA4DD: data_out = 8'h81;
                    16'hA4DE: data_out = 8'h82;
                    16'hA4DF: data_out = 8'h83;
                    16'hA4E0: data_out = 8'h84;
                    16'hA4E1: data_out = 8'h85;
                    16'hA4E2: data_out = 8'h86;
                    16'hA4E3: data_out = 8'h87;
                    16'hA4E4: data_out = 8'h88;
                    16'hA4E5: data_out = 8'h89;
                    16'hA4E6: data_out = 8'h8A;
                    16'hA4E7: data_out = 8'h8B;
                    16'hA4E8: data_out = 8'h8C;
                    16'hA4E9: data_out = 8'h8D;
                    16'hA4EA: data_out = 8'h8E;
                    16'hA4EB: data_out = 8'h8F;
                    16'hA4EC: data_out = 8'h90;
                    16'hA4ED: data_out = 8'h91;
                    16'hA4EE: data_out = 8'h92;
                    16'hA4EF: data_out = 8'h93;
                    16'hA4F0: data_out = 8'h94;
                    16'hA4F1: data_out = 8'h95;
                    16'hA4F2: data_out = 8'h96;
                    16'hA4F3: data_out = 8'h97;
                    16'hA4F4: data_out = 8'h98;
                    16'hA4F5: data_out = 8'h99;
                    16'hA4F6: data_out = 8'h9A;
                    16'hA4F7: data_out = 8'h9B;
                    16'hA4F8: data_out = 8'h9C;
                    16'hA4F9: data_out = 8'h9D;
                    16'hA4FA: data_out = 8'h9E;
                    16'hA4FB: data_out = 8'h9F;
                    16'hA4FC: data_out = 8'hA0;
                    16'hA4FD: data_out = 8'hA1;
                    16'hA4FE: data_out = 8'hA2;
                    16'hA4FF: data_out = 8'hA3;
                    16'hA500: data_out = 8'hA5;
                    16'hA501: data_out = 8'hA4;
                    16'hA502: data_out = 8'hA3;
                    16'hA503: data_out = 8'hA2;
                    16'hA504: data_out = 8'hA1;
                    16'hA505: data_out = 8'hA0;
                    16'hA506: data_out = 8'h9F;
                    16'hA507: data_out = 8'h9E;
                    16'hA508: data_out = 8'h9D;
                    16'hA509: data_out = 8'h9C;
                    16'hA50A: data_out = 8'h9B;
                    16'hA50B: data_out = 8'h9A;
                    16'hA50C: data_out = 8'h99;
                    16'hA50D: data_out = 8'h98;
                    16'hA50E: data_out = 8'h97;
                    16'hA50F: data_out = 8'h96;
                    16'hA510: data_out = 8'h95;
                    16'hA511: data_out = 8'h94;
                    16'hA512: data_out = 8'h93;
                    16'hA513: data_out = 8'h92;
                    16'hA514: data_out = 8'h91;
                    16'hA515: data_out = 8'h90;
                    16'hA516: data_out = 8'h8F;
                    16'hA517: data_out = 8'h8E;
                    16'hA518: data_out = 8'h8D;
                    16'hA519: data_out = 8'h8C;
                    16'hA51A: data_out = 8'h8B;
                    16'hA51B: data_out = 8'h8A;
                    16'hA51C: data_out = 8'h89;
                    16'hA51D: data_out = 8'h88;
                    16'hA51E: data_out = 8'h87;
                    16'hA51F: data_out = 8'h86;
                    16'hA520: data_out = 8'h85;
                    16'hA521: data_out = 8'h84;
                    16'hA522: data_out = 8'h83;
                    16'hA523: data_out = 8'h82;
                    16'hA524: data_out = 8'h81;
                    16'hA525: data_out = 8'h0;
                    16'hA526: data_out = 8'h1;
                    16'hA527: data_out = 8'h2;
                    16'hA528: data_out = 8'h3;
                    16'hA529: data_out = 8'h4;
                    16'hA52A: data_out = 8'h5;
                    16'hA52B: data_out = 8'h6;
                    16'hA52C: data_out = 8'h7;
                    16'hA52D: data_out = 8'h8;
                    16'hA52E: data_out = 8'h9;
                    16'hA52F: data_out = 8'hA;
                    16'hA530: data_out = 8'hB;
                    16'hA531: data_out = 8'hC;
                    16'hA532: data_out = 8'hD;
                    16'hA533: data_out = 8'hE;
                    16'hA534: data_out = 8'hF;
                    16'hA535: data_out = 8'h10;
                    16'hA536: data_out = 8'h11;
                    16'hA537: data_out = 8'h12;
                    16'hA538: data_out = 8'h13;
                    16'hA539: data_out = 8'h14;
                    16'hA53A: data_out = 8'h15;
                    16'hA53B: data_out = 8'h16;
                    16'hA53C: data_out = 8'h17;
                    16'hA53D: data_out = 8'h18;
                    16'hA53E: data_out = 8'h19;
                    16'hA53F: data_out = 8'h1A;
                    16'hA540: data_out = 8'h1B;
                    16'hA541: data_out = 8'h1C;
                    16'hA542: data_out = 8'h1D;
                    16'hA543: data_out = 8'h1E;
                    16'hA544: data_out = 8'h1F;
                    16'hA545: data_out = 8'h20;
                    16'hA546: data_out = 8'h21;
                    16'hA547: data_out = 8'h22;
                    16'hA548: data_out = 8'h23;
                    16'hA549: data_out = 8'h24;
                    16'hA54A: data_out = 8'h25;
                    16'hA54B: data_out = 8'h26;
                    16'hA54C: data_out = 8'h27;
                    16'hA54D: data_out = 8'h28;
                    16'hA54E: data_out = 8'h29;
                    16'hA54F: data_out = 8'h2A;
                    16'hA550: data_out = 8'h2B;
                    16'hA551: data_out = 8'h2C;
                    16'hA552: data_out = 8'h2D;
                    16'hA553: data_out = 8'h2E;
                    16'hA554: data_out = 8'h2F;
                    16'hA555: data_out = 8'h30;
                    16'hA556: data_out = 8'h31;
                    16'hA557: data_out = 8'h32;
                    16'hA558: data_out = 8'h33;
                    16'hA559: data_out = 8'h34;
                    16'hA55A: data_out = 8'h35;
                    16'hA55B: data_out = 8'h36;
                    16'hA55C: data_out = 8'h37;
                    16'hA55D: data_out = 8'h38;
                    16'hA55E: data_out = 8'h39;
                    16'hA55F: data_out = 8'h3A;
                    16'hA560: data_out = 8'h3B;
                    16'hA561: data_out = 8'h3C;
                    16'hA562: data_out = 8'h3D;
                    16'hA563: data_out = 8'h3E;
                    16'hA564: data_out = 8'h3F;
                    16'hA565: data_out = 8'h40;
                    16'hA566: data_out = 8'h41;
                    16'hA567: data_out = 8'h42;
                    16'hA568: data_out = 8'h43;
                    16'hA569: data_out = 8'h44;
                    16'hA56A: data_out = 8'h45;
                    16'hA56B: data_out = 8'h46;
                    16'hA56C: data_out = 8'h47;
                    16'hA56D: data_out = 8'h48;
                    16'hA56E: data_out = 8'h49;
                    16'hA56F: data_out = 8'h4A;
                    16'hA570: data_out = 8'h4B;
                    16'hA571: data_out = 8'h4C;
                    16'hA572: data_out = 8'h4D;
                    16'hA573: data_out = 8'h4E;
                    16'hA574: data_out = 8'h4F;
                    16'hA575: data_out = 8'h50;
                    16'hA576: data_out = 8'h51;
                    16'hA577: data_out = 8'h52;
                    16'hA578: data_out = 8'h53;
                    16'hA579: data_out = 8'h54;
                    16'hA57A: data_out = 8'h55;
                    16'hA57B: data_out = 8'h56;
                    16'hA57C: data_out = 8'h57;
                    16'hA57D: data_out = 8'h58;
                    16'hA57E: data_out = 8'h59;
                    16'hA57F: data_out = 8'h5A;
                    16'hA580: data_out = 8'hA5;
                    16'hA581: data_out = 8'hA6;
                    16'hA582: data_out = 8'hA7;
                    16'hA583: data_out = 8'hA8;
                    16'hA584: data_out = 8'hA9;
                    16'hA585: data_out = 8'hAA;
                    16'hA586: data_out = 8'hAB;
                    16'hA587: data_out = 8'hAC;
                    16'hA588: data_out = 8'hAD;
                    16'hA589: data_out = 8'hAE;
                    16'hA58A: data_out = 8'hAF;
                    16'hA58B: data_out = 8'hB0;
                    16'hA58C: data_out = 8'hB1;
                    16'hA58D: data_out = 8'hB2;
                    16'hA58E: data_out = 8'hB3;
                    16'hA58F: data_out = 8'hB4;
                    16'hA590: data_out = 8'hB5;
                    16'hA591: data_out = 8'hB6;
                    16'hA592: data_out = 8'hB7;
                    16'hA593: data_out = 8'hB8;
                    16'hA594: data_out = 8'hB9;
                    16'hA595: data_out = 8'hBA;
                    16'hA596: data_out = 8'hBB;
                    16'hA597: data_out = 8'hBC;
                    16'hA598: data_out = 8'hBD;
                    16'hA599: data_out = 8'hBE;
                    16'hA59A: data_out = 8'hBF;
                    16'hA59B: data_out = 8'hC0;
                    16'hA59C: data_out = 8'hC1;
                    16'hA59D: data_out = 8'hC2;
                    16'hA59E: data_out = 8'hC3;
                    16'hA59F: data_out = 8'hC4;
                    16'hA5A0: data_out = 8'hC5;
                    16'hA5A1: data_out = 8'hC6;
                    16'hA5A2: data_out = 8'hC7;
                    16'hA5A3: data_out = 8'hC8;
                    16'hA5A4: data_out = 8'hC9;
                    16'hA5A5: data_out = 8'hCA;
                    16'hA5A6: data_out = 8'hCB;
                    16'hA5A7: data_out = 8'hCC;
                    16'hA5A8: data_out = 8'hCD;
                    16'hA5A9: data_out = 8'hCE;
                    16'hA5AA: data_out = 8'hCF;
                    16'hA5AB: data_out = 8'hD0;
                    16'hA5AC: data_out = 8'hD1;
                    16'hA5AD: data_out = 8'hD2;
                    16'hA5AE: data_out = 8'hD3;
                    16'hA5AF: data_out = 8'hD4;
                    16'hA5B0: data_out = 8'hD5;
                    16'hA5B1: data_out = 8'hD6;
                    16'hA5B2: data_out = 8'hD7;
                    16'hA5B3: data_out = 8'hD8;
                    16'hA5B4: data_out = 8'hD9;
                    16'hA5B5: data_out = 8'hDA;
                    16'hA5B6: data_out = 8'hDB;
                    16'hA5B7: data_out = 8'hDC;
                    16'hA5B8: data_out = 8'hDD;
                    16'hA5B9: data_out = 8'hDE;
                    16'hA5BA: data_out = 8'hDF;
                    16'hA5BB: data_out = 8'hE0;
                    16'hA5BC: data_out = 8'hE1;
                    16'hA5BD: data_out = 8'hE2;
                    16'hA5BE: data_out = 8'hE3;
                    16'hA5BF: data_out = 8'hE4;
                    16'hA5C0: data_out = 8'hE5;
                    16'hA5C1: data_out = 8'hE6;
                    16'hA5C2: data_out = 8'hE7;
                    16'hA5C3: data_out = 8'hE8;
                    16'hA5C4: data_out = 8'hE9;
                    16'hA5C5: data_out = 8'hEA;
                    16'hA5C6: data_out = 8'hEB;
                    16'hA5C7: data_out = 8'hEC;
                    16'hA5C8: data_out = 8'hED;
                    16'hA5C9: data_out = 8'hEE;
                    16'hA5CA: data_out = 8'hEF;
                    16'hA5CB: data_out = 8'hF0;
                    16'hA5CC: data_out = 8'hF1;
                    16'hA5CD: data_out = 8'hF2;
                    16'hA5CE: data_out = 8'hF3;
                    16'hA5CF: data_out = 8'hF4;
                    16'hA5D0: data_out = 8'hF5;
                    16'hA5D1: data_out = 8'hF6;
                    16'hA5D2: data_out = 8'hF7;
                    16'hA5D3: data_out = 8'hF8;
                    16'hA5D4: data_out = 8'hF9;
                    16'hA5D5: data_out = 8'hFA;
                    16'hA5D6: data_out = 8'hFB;
                    16'hA5D7: data_out = 8'hFC;
                    16'hA5D8: data_out = 8'hFD;
                    16'hA5D9: data_out = 8'hFE;
                    16'hA5DA: data_out = 8'hFF;
                    16'hA5DB: data_out = 8'h80;
                    16'hA5DC: data_out = 8'h81;
                    16'hA5DD: data_out = 8'h82;
                    16'hA5DE: data_out = 8'h83;
                    16'hA5DF: data_out = 8'h84;
                    16'hA5E0: data_out = 8'h85;
                    16'hA5E1: data_out = 8'h86;
                    16'hA5E2: data_out = 8'h87;
                    16'hA5E3: data_out = 8'h88;
                    16'hA5E4: data_out = 8'h89;
                    16'hA5E5: data_out = 8'h8A;
                    16'hA5E6: data_out = 8'h8B;
                    16'hA5E7: data_out = 8'h8C;
                    16'hA5E8: data_out = 8'h8D;
                    16'hA5E9: data_out = 8'h8E;
                    16'hA5EA: data_out = 8'h8F;
                    16'hA5EB: data_out = 8'h90;
                    16'hA5EC: data_out = 8'h91;
                    16'hA5ED: data_out = 8'h92;
                    16'hA5EE: data_out = 8'h93;
                    16'hA5EF: data_out = 8'h94;
                    16'hA5F0: data_out = 8'h95;
                    16'hA5F1: data_out = 8'h96;
                    16'hA5F2: data_out = 8'h97;
                    16'hA5F3: data_out = 8'h98;
                    16'hA5F4: data_out = 8'h99;
                    16'hA5F5: data_out = 8'h9A;
                    16'hA5F6: data_out = 8'h9B;
                    16'hA5F7: data_out = 8'h9C;
                    16'hA5F8: data_out = 8'h9D;
                    16'hA5F9: data_out = 8'h9E;
                    16'hA5FA: data_out = 8'h9F;
                    16'hA5FB: data_out = 8'hA0;
                    16'hA5FC: data_out = 8'hA1;
                    16'hA5FD: data_out = 8'hA2;
                    16'hA5FE: data_out = 8'hA3;
                    16'hA5FF: data_out = 8'hA4;
                    16'hA600: data_out = 8'hA6;
                    16'hA601: data_out = 8'hA5;
                    16'hA602: data_out = 8'hA4;
                    16'hA603: data_out = 8'hA3;
                    16'hA604: data_out = 8'hA2;
                    16'hA605: data_out = 8'hA1;
                    16'hA606: data_out = 8'hA0;
                    16'hA607: data_out = 8'h9F;
                    16'hA608: data_out = 8'h9E;
                    16'hA609: data_out = 8'h9D;
                    16'hA60A: data_out = 8'h9C;
                    16'hA60B: data_out = 8'h9B;
                    16'hA60C: data_out = 8'h9A;
                    16'hA60D: data_out = 8'h99;
                    16'hA60E: data_out = 8'h98;
                    16'hA60F: data_out = 8'h97;
                    16'hA610: data_out = 8'h96;
                    16'hA611: data_out = 8'h95;
                    16'hA612: data_out = 8'h94;
                    16'hA613: data_out = 8'h93;
                    16'hA614: data_out = 8'h92;
                    16'hA615: data_out = 8'h91;
                    16'hA616: data_out = 8'h90;
                    16'hA617: data_out = 8'h8F;
                    16'hA618: data_out = 8'h8E;
                    16'hA619: data_out = 8'h8D;
                    16'hA61A: data_out = 8'h8C;
                    16'hA61B: data_out = 8'h8B;
                    16'hA61C: data_out = 8'h8A;
                    16'hA61D: data_out = 8'h89;
                    16'hA61E: data_out = 8'h88;
                    16'hA61F: data_out = 8'h87;
                    16'hA620: data_out = 8'h86;
                    16'hA621: data_out = 8'h85;
                    16'hA622: data_out = 8'h84;
                    16'hA623: data_out = 8'h83;
                    16'hA624: data_out = 8'h82;
                    16'hA625: data_out = 8'h81;
                    16'hA626: data_out = 8'h0;
                    16'hA627: data_out = 8'h1;
                    16'hA628: data_out = 8'h2;
                    16'hA629: data_out = 8'h3;
                    16'hA62A: data_out = 8'h4;
                    16'hA62B: data_out = 8'h5;
                    16'hA62C: data_out = 8'h6;
                    16'hA62D: data_out = 8'h7;
                    16'hA62E: data_out = 8'h8;
                    16'hA62F: data_out = 8'h9;
                    16'hA630: data_out = 8'hA;
                    16'hA631: data_out = 8'hB;
                    16'hA632: data_out = 8'hC;
                    16'hA633: data_out = 8'hD;
                    16'hA634: data_out = 8'hE;
                    16'hA635: data_out = 8'hF;
                    16'hA636: data_out = 8'h10;
                    16'hA637: data_out = 8'h11;
                    16'hA638: data_out = 8'h12;
                    16'hA639: data_out = 8'h13;
                    16'hA63A: data_out = 8'h14;
                    16'hA63B: data_out = 8'h15;
                    16'hA63C: data_out = 8'h16;
                    16'hA63D: data_out = 8'h17;
                    16'hA63E: data_out = 8'h18;
                    16'hA63F: data_out = 8'h19;
                    16'hA640: data_out = 8'h1A;
                    16'hA641: data_out = 8'h1B;
                    16'hA642: data_out = 8'h1C;
                    16'hA643: data_out = 8'h1D;
                    16'hA644: data_out = 8'h1E;
                    16'hA645: data_out = 8'h1F;
                    16'hA646: data_out = 8'h20;
                    16'hA647: data_out = 8'h21;
                    16'hA648: data_out = 8'h22;
                    16'hA649: data_out = 8'h23;
                    16'hA64A: data_out = 8'h24;
                    16'hA64B: data_out = 8'h25;
                    16'hA64C: data_out = 8'h26;
                    16'hA64D: data_out = 8'h27;
                    16'hA64E: data_out = 8'h28;
                    16'hA64F: data_out = 8'h29;
                    16'hA650: data_out = 8'h2A;
                    16'hA651: data_out = 8'h2B;
                    16'hA652: data_out = 8'h2C;
                    16'hA653: data_out = 8'h2D;
                    16'hA654: data_out = 8'h2E;
                    16'hA655: data_out = 8'h2F;
                    16'hA656: data_out = 8'h30;
                    16'hA657: data_out = 8'h31;
                    16'hA658: data_out = 8'h32;
                    16'hA659: data_out = 8'h33;
                    16'hA65A: data_out = 8'h34;
                    16'hA65B: data_out = 8'h35;
                    16'hA65C: data_out = 8'h36;
                    16'hA65D: data_out = 8'h37;
                    16'hA65E: data_out = 8'h38;
                    16'hA65F: data_out = 8'h39;
                    16'hA660: data_out = 8'h3A;
                    16'hA661: data_out = 8'h3B;
                    16'hA662: data_out = 8'h3C;
                    16'hA663: data_out = 8'h3D;
                    16'hA664: data_out = 8'h3E;
                    16'hA665: data_out = 8'h3F;
                    16'hA666: data_out = 8'h40;
                    16'hA667: data_out = 8'h41;
                    16'hA668: data_out = 8'h42;
                    16'hA669: data_out = 8'h43;
                    16'hA66A: data_out = 8'h44;
                    16'hA66B: data_out = 8'h45;
                    16'hA66C: data_out = 8'h46;
                    16'hA66D: data_out = 8'h47;
                    16'hA66E: data_out = 8'h48;
                    16'hA66F: data_out = 8'h49;
                    16'hA670: data_out = 8'h4A;
                    16'hA671: data_out = 8'h4B;
                    16'hA672: data_out = 8'h4C;
                    16'hA673: data_out = 8'h4D;
                    16'hA674: data_out = 8'h4E;
                    16'hA675: data_out = 8'h4F;
                    16'hA676: data_out = 8'h50;
                    16'hA677: data_out = 8'h51;
                    16'hA678: data_out = 8'h52;
                    16'hA679: data_out = 8'h53;
                    16'hA67A: data_out = 8'h54;
                    16'hA67B: data_out = 8'h55;
                    16'hA67C: data_out = 8'h56;
                    16'hA67D: data_out = 8'h57;
                    16'hA67E: data_out = 8'h58;
                    16'hA67F: data_out = 8'h59;
                    16'hA680: data_out = 8'hA6;
                    16'hA681: data_out = 8'hA7;
                    16'hA682: data_out = 8'hA8;
                    16'hA683: data_out = 8'hA9;
                    16'hA684: data_out = 8'hAA;
                    16'hA685: data_out = 8'hAB;
                    16'hA686: data_out = 8'hAC;
                    16'hA687: data_out = 8'hAD;
                    16'hA688: data_out = 8'hAE;
                    16'hA689: data_out = 8'hAF;
                    16'hA68A: data_out = 8'hB0;
                    16'hA68B: data_out = 8'hB1;
                    16'hA68C: data_out = 8'hB2;
                    16'hA68D: data_out = 8'hB3;
                    16'hA68E: data_out = 8'hB4;
                    16'hA68F: data_out = 8'hB5;
                    16'hA690: data_out = 8'hB6;
                    16'hA691: data_out = 8'hB7;
                    16'hA692: data_out = 8'hB8;
                    16'hA693: data_out = 8'hB9;
                    16'hA694: data_out = 8'hBA;
                    16'hA695: data_out = 8'hBB;
                    16'hA696: data_out = 8'hBC;
                    16'hA697: data_out = 8'hBD;
                    16'hA698: data_out = 8'hBE;
                    16'hA699: data_out = 8'hBF;
                    16'hA69A: data_out = 8'hC0;
                    16'hA69B: data_out = 8'hC1;
                    16'hA69C: data_out = 8'hC2;
                    16'hA69D: data_out = 8'hC3;
                    16'hA69E: data_out = 8'hC4;
                    16'hA69F: data_out = 8'hC5;
                    16'hA6A0: data_out = 8'hC6;
                    16'hA6A1: data_out = 8'hC7;
                    16'hA6A2: data_out = 8'hC8;
                    16'hA6A3: data_out = 8'hC9;
                    16'hA6A4: data_out = 8'hCA;
                    16'hA6A5: data_out = 8'hCB;
                    16'hA6A6: data_out = 8'hCC;
                    16'hA6A7: data_out = 8'hCD;
                    16'hA6A8: data_out = 8'hCE;
                    16'hA6A9: data_out = 8'hCF;
                    16'hA6AA: data_out = 8'hD0;
                    16'hA6AB: data_out = 8'hD1;
                    16'hA6AC: data_out = 8'hD2;
                    16'hA6AD: data_out = 8'hD3;
                    16'hA6AE: data_out = 8'hD4;
                    16'hA6AF: data_out = 8'hD5;
                    16'hA6B0: data_out = 8'hD6;
                    16'hA6B1: data_out = 8'hD7;
                    16'hA6B2: data_out = 8'hD8;
                    16'hA6B3: data_out = 8'hD9;
                    16'hA6B4: data_out = 8'hDA;
                    16'hA6B5: data_out = 8'hDB;
                    16'hA6B6: data_out = 8'hDC;
                    16'hA6B7: data_out = 8'hDD;
                    16'hA6B8: data_out = 8'hDE;
                    16'hA6B9: data_out = 8'hDF;
                    16'hA6BA: data_out = 8'hE0;
                    16'hA6BB: data_out = 8'hE1;
                    16'hA6BC: data_out = 8'hE2;
                    16'hA6BD: data_out = 8'hE3;
                    16'hA6BE: data_out = 8'hE4;
                    16'hA6BF: data_out = 8'hE5;
                    16'hA6C0: data_out = 8'hE6;
                    16'hA6C1: data_out = 8'hE7;
                    16'hA6C2: data_out = 8'hE8;
                    16'hA6C3: data_out = 8'hE9;
                    16'hA6C4: data_out = 8'hEA;
                    16'hA6C5: data_out = 8'hEB;
                    16'hA6C6: data_out = 8'hEC;
                    16'hA6C7: data_out = 8'hED;
                    16'hA6C8: data_out = 8'hEE;
                    16'hA6C9: data_out = 8'hEF;
                    16'hA6CA: data_out = 8'hF0;
                    16'hA6CB: data_out = 8'hF1;
                    16'hA6CC: data_out = 8'hF2;
                    16'hA6CD: data_out = 8'hF3;
                    16'hA6CE: data_out = 8'hF4;
                    16'hA6CF: data_out = 8'hF5;
                    16'hA6D0: data_out = 8'hF6;
                    16'hA6D1: data_out = 8'hF7;
                    16'hA6D2: data_out = 8'hF8;
                    16'hA6D3: data_out = 8'hF9;
                    16'hA6D4: data_out = 8'hFA;
                    16'hA6D5: data_out = 8'hFB;
                    16'hA6D6: data_out = 8'hFC;
                    16'hA6D7: data_out = 8'hFD;
                    16'hA6D8: data_out = 8'hFE;
                    16'hA6D9: data_out = 8'hFF;
                    16'hA6DA: data_out = 8'h80;
                    16'hA6DB: data_out = 8'h81;
                    16'hA6DC: data_out = 8'h82;
                    16'hA6DD: data_out = 8'h83;
                    16'hA6DE: data_out = 8'h84;
                    16'hA6DF: data_out = 8'h85;
                    16'hA6E0: data_out = 8'h86;
                    16'hA6E1: data_out = 8'h87;
                    16'hA6E2: data_out = 8'h88;
                    16'hA6E3: data_out = 8'h89;
                    16'hA6E4: data_out = 8'h8A;
                    16'hA6E5: data_out = 8'h8B;
                    16'hA6E6: data_out = 8'h8C;
                    16'hA6E7: data_out = 8'h8D;
                    16'hA6E8: data_out = 8'h8E;
                    16'hA6E9: data_out = 8'h8F;
                    16'hA6EA: data_out = 8'h90;
                    16'hA6EB: data_out = 8'h91;
                    16'hA6EC: data_out = 8'h92;
                    16'hA6ED: data_out = 8'h93;
                    16'hA6EE: data_out = 8'h94;
                    16'hA6EF: data_out = 8'h95;
                    16'hA6F0: data_out = 8'h96;
                    16'hA6F1: data_out = 8'h97;
                    16'hA6F2: data_out = 8'h98;
                    16'hA6F3: data_out = 8'h99;
                    16'hA6F4: data_out = 8'h9A;
                    16'hA6F5: data_out = 8'h9B;
                    16'hA6F6: data_out = 8'h9C;
                    16'hA6F7: data_out = 8'h9D;
                    16'hA6F8: data_out = 8'h9E;
                    16'hA6F9: data_out = 8'h9F;
                    16'hA6FA: data_out = 8'hA0;
                    16'hA6FB: data_out = 8'hA1;
                    16'hA6FC: data_out = 8'hA2;
                    16'hA6FD: data_out = 8'hA3;
                    16'hA6FE: data_out = 8'hA4;
                    16'hA6FF: data_out = 8'hA5;
                    16'hA700: data_out = 8'hA7;
                    16'hA701: data_out = 8'hA6;
                    16'hA702: data_out = 8'hA5;
                    16'hA703: data_out = 8'hA4;
                    16'hA704: data_out = 8'hA3;
                    16'hA705: data_out = 8'hA2;
                    16'hA706: data_out = 8'hA1;
                    16'hA707: data_out = 8'hA0;
                    16'hA708: data_out = 8'h9F;
                    16'hA709: data_out = 8'h9E;
                    16'hA70A: data_out = 8'h9D;
                    16'hA70B: data_out = 8'h9C;
                    16'hA70C: data_out = 8'h9B;
                    16'hA70D: data_out = 8'h9A;
                    16'hA70E: data_out = 8'h99;
                    16'hA70F: data_out = 8'h98;
                    16'hA710: data_out = 8'h97;
                    16'hA711: data_out = 8'h96;
                    16'hA712: data_out = 8'h95;
                    16'hA713: data_out = 8'h94;
                    16'hA714: data_out = 8'h93;
                    16'hA715: data_out = 8'h92;
                    16'hA716: data_out = 8'h91;
                    16'hA717: data_out = 8'h90;
                    16'hA718: data_out = 8'h8F;
                    16'hA719: data_out = 8'h8E;
                    16'hA71A: data_out = 8'h8D;
                    16'hA71B: data_out = 8'h8C;
                    16'hA71C: data_out = 8'h8B;
                    16'hA71D: data_out = 8'h8A;
                    16'hA71E: data_out = 8'h89;
                    16'hA71F: data_out = 8'h88;
                    16'hA720: data_out = 8'h87;
                    16'hA721: data_out = 8'h86;
                    16'hA722: data_out = 8'h85;
                    16'hA723: data_out = 8'h84;
                    16'hA724: data_out = 8'h83;
                    16'hA725: data_out = 8'h82;
                    16'hA726: data_out = 8'h81;
                    16'hA727: data_out = 8'h0;
                    16'hA728: data_out = 8'h1;
                    16'hA729: data_out = 8'h2;
                    16'hA72A: data_out = 8'h3;
                    16'hA72B: data_out = 8'h4;
                    16'hA72C: data_out = 8'h5;
                    16'hA72D: data_out = 8'h6;
                    16'hA72E: data_out = 8'h7;
                    16'hA72F: data_out = 8'h8;
                    16'hA730: data_out = 8'h9;
                    16'hA731: data_out = 8'hA;
                    16'hA732: data_out = 8'hB;
                    16'hA733: data_out = 8'hC;
                    16'hA734: data_out = 8'hD;
                    16'hA735: data_out = 8'hE;
                    16'hA736: data_out = 8'hF;
                    16'hA737: data_out = 8'h10;
                    16'hA738: data_out = 8'h11;
                    16'hA739: data_out = 8'h12;
                    16'hA73A: data_out = 8'h13;
                    16'hA73B: data_out = 8'h14;
                    16'hA73C: data_out = 8'h15;
                    16'hA73D: data_out = 8'h16;
                    16'hA73E: data_out = 8'h17;
                    16'hA73F: data_out = 8'h18;
                    16'hA740: data_out = 8'h19;
                    16'hA741: data_out = 8'h1A;
                    16'hA742: data_out = 8'h1B;
                    16'hA743: data_out = 8'h1C;
                    16'hA744: data_out = 8'h1D;
                    16'hA745: data_out = 8'h1E;
                    16'hA746: data_out = 8'h1F;
                    16'hA747: data_out = 8'h20;
                    16'hA748: data_out = 8'h21;
                    16'hA749: data_out = 8'h22;
                    16'hA74A: data_out = 8'h23;
                    16'hA74B: data_out = 8'h24;
                    16'hA74C: data_out = 8'h25;
                    16'hA74D: data_out = 8'h26;
                    16'hA74E: data_out = 8'h27;
                    16'hA74F: data_out = 8'h28;
                    16'hA750: data_out = 8'h29;
                    16'hA751: data_out = 8'h2A;
                    16'hA752: data_out = 8'h2B;
                    16'hA753: data_out = 8'h2C;
                    16'hA754: data_out = 8'h2D;
                    16'hA755: data_out = 8'h2E;
                    16'hA756: data_out = 8'h2F;
                    16'hA757: data_out = 8'h30;
                    16'hA758: data_out = 8'h31;
                    16'hA759: data_out = 8'h32;
                    16'hA75A: data_out = 8'h33;
                    16'hA75B: data_out = 8'h34;
                    16'hA75C: data_out = 8'h35;
                    16'hA75D: data_out = 8'h36;
                    16'hA75E: data_out = 8'h37;
                    16'hA75F: data_out = 8'h38;
                    16'hA760: data_out = 8'h39;
                    16'hA761: data_out = 8'h3A;
                    16'hA762: data_out = 8'h3B;
                    16'hA763: data_out = 8'h3C;
                    16'hA764: data_out = 8'h3D;
                    16'hA765: data_out = 8'h3E;
                    16'hA766: data_out = 8'h3F;
                    16'hA767: data_out = 8'h40;
                    16'hA768: data_out = 8'h41;
                    16'hA769: data_out = 8'h42;
                    16'hA76A: data_out = 8'h43;
                    16'hA76B: data_out = 8'h44;
                    16'hA76C: data_out = 8'h45;
                    16'hA76D: data_out = 8'h46;
                    16'hA76E: data_out = 8'h47;
                    16'hA76F: data_out = 8'h48;
                    16'hA770: data_out = 8'h49;
                    16'hA771: data_out = 8'h4A;
                    16'hA772: data_out = 8'h4B;
                    16'hA773: data_out = 8'h4C;
                    16'hA774: data_out = 8'h4D;
                    16'hA775: data_out = 8'h4E;
                    16'hA776: data_out = 8'h4F;
                    16'hA777: data_out = 8'h50;
                    16'hA778: data_out = 8'h51;
                    16'hA779: data_out = 8'h52;
                    16'hA77A: data_out = 8'h53;
                    16'hA77B: data_out = 8'h54;
                    16'hA77C: data_out = 8'h55;
                    16'hA77D: data_out = 8'h56;
                    16'hA77E: data_out = 8'h57;
                    16'hA77F: data_out = 8'h58;
                    16'hA780: data_out = 8'hA7;
                    16'hA781: data_out = 8'hA8;
                    16'hA782: data_out = 8'hA9;
                    16'hA783: data_out = 8'hAA;
                    16'hA784: data_out = 8'hAB;
                    16'hA785: data_out = 8'hAC;
                    16'hA786: data_out = 8'hAD;
                    16'hA787: data_out = 8'hAE;
                    16'hA788: data_out = 8'hAF;
                    16'hA789: data_out = 8'hB0;
                    16'hA78A: data_out = 8'hB1;
                    16'hA78B: data_out = 8'hB2;
                    16'hA78C: data_out = 8'hB3;
                    16'hA78D: data_out = 8'hB4;
                    16'hA78E: data_out = 8'hB5;
                    16'hA78F: data_out = 8'hB6;
                    16'hA790: data_out = 8'hB7;
                    16'hA791: data_out = 8'hB8;
                    16'hA792: data_out = 8'hB9;
                    16'hA793: data_out = 8'hBA;
                    16'hA794: data_out = 8'hBB;
                    16'hA795: data_out = 8'hBC;
                    16'hA796: data_out = 8'hBD;
                    16'hA797: data_out = 8'hBE;
                    16'hA798: data_out = 8'hBF;
                    16'hA799: data_out = 8'hC0;
                    16'hA79A: data_out = 8'hC1;
                    16'hA79B: data_out = 8'hC2;
                    16'hA79C: data_out = 8'hC3;
                    16'hA79D: data_out = 8'hC4;
                    16'hA79E: data_out = 8'hC5;
                    16'hA79F: data_out = 8'hC6;
                    16'hA7A0: data_out = 8'hC7;
                    16'hA7A1: data_out = 8'hC8;
                    16'hA7A2: data_out = 8'hC9;
                    16'hA7A3: data_out = 8'hCA;
                    16'hA7A4: data_out = 8'hCB;
                    16'hA7A5: data_out = 8'hCC;
                    16'hA7A6: data_out = 8'hCD;
                    16'hA7A7: data_out = 8'hCE;
                    16'hA7A8: data_out = 8'hCF;
                    16'hA7A9: data_out = 8'hD0;
                    16'hA7AA: data_out = 8'hD1;
                    16'hA7AB: data_out = 8'hD2;
                    16'hA7AC: data_out = 8'hD3;
                    16'hA7AD: data_out = 8'hD4;
                    16'hA7AE: data_out = 8'hD5;
                    16'hA7AF: data_out = 8'hD6;
                    16'hA7B0: data_out = 8'hD7;
                    16'hA7B1: data_out = 8'hD8;
                    16'hA7B2: data_out = 8'hD9;
                    16'hA7B3: data_out = 8'hDA;
                    16'hA7B4: data_out = 8'hDB;
                    16'hA7B5: data_out = 8'hDC;
                    16'hA7B6: data_out = 8'hDD;
                    16'hA7B7: data_out = 8'hDE;
                    16'hA7B8: data_out = 8'hDF;
                    16'hA7B9: data_out = 8'hE0;
                    16'hA7BA: data_out = 8'hE1;
                    16'hA7BB: data_out = 8'hE2;
                    16'hA7BC: data_out = 8'hE3;
                    16'hA7BD: data_out = 8'hE4;
                    16'hA7BE: data_out = 8'hE5;
                    16'hA7BF: data_out = 8'hE6;
                    16'hA7C0: data_out = 8'hE7;
                    16'hA7C1: data_out = 8'hE8;
                    16'hA7C2: data_out = 8'hE9;
                    16'hA7C3: data_out = 8'hEA;
                    16'hA7C4: data_out = 8'hEB;
                    16'hA7C5: data_out = 8'hEC;
                    16'hA7C6: data_out = 8'hED;
                    16'hA7C7: data_out = 8'hEE;
                    16'hA7C8: data_out = 8'hEF;
                    16'hA7C9: data_out = 8'hF0;
                    16'hA7CA: data_out = 8'hF1;
                    16'hA7CB: data_out = 8'hF2;
                    16'hA7CC: data_out = 8'hF3;
                    16'hA7CD: data_out = 8'hF4;
                    16'hA7CE: data_out = 8'hF5;
                    16'hA7CF: data_out = 8'hF6;
                    16'hA7D0: data_out = 8'hF7;
                    16'hA7D1: data_out = 8'hF8;
                    16'hA7D2: data_out = 8'hF9;
                    16'hA7D3: data_out = 8'hFA;
                    16'hA7D4: data_out = 8'hFB;
                    16'hA7D5: data_out = 8'hFC;
                    16'hA7D6: data_out = 8'hFD;
                    16'hA7D7: data_out = 8'hFE;
                    16'hA7D8: data_out = 8'hFF;
                    16'hA7D9: data_out = 8'h80;
                    16'hA7DA: data_out = 8'h81;
                    16'hA7DB: data_out = 8'h82;
                    16'hA7DC: data_out = 8'h83;
                    16'hA7DD: data_out = 8'h84;
                    16'hA7DE: data_out = 8'h85;
                    16'hA7DF: data_out = 8'h86;
                    16'hA7E0: data_out = 8'h87;
                    16'hA7E1: data_out = 8'h88;
                    16'hA7E2: data_out = 8'h89;
                    16'hA7E3: data_out = 8'h8A;
                    16'hA7E4: data_out = 8'h8B;
                    16'hA7E5: data_out = 8'h8C;
                    16'hA7E6: data_out = 8'h8D;
                    16'hA7E7: data_out = 8'h8E;
                    16'hA7E8: data_out = 8'h8F;
                    16'hA7E9: data_out = 8'h90;
                    16'hA7EA: data_out = 8'h91;
                    16'hA7EB: data_out = 8'h92;
                    16'hA7EC: data_out = 8'h93;
                    16'hA7ED: data_out = 8'h94;
                    16'hA7EE: data_out = 8'h95;
                    16'hA7EF: data_out = 8'h96;
                    16'hA7F0: data_out = 8'h97;
                    16'hA7F1: data_out = 8'h98;
                    16'hA7F2: data_out = 8'h99;
                    16'hA7F3: data_out = 8'h9A;
                    16'hA7F4: data_out = 8'h9B;
                    16'hA7F5: data_out = 8'h9C;
                    16'hA7F6: data_out = 8'h9D;
                    16'hA7F7: data_out = 8'h9E;
                    16'hA7F8: data_out = 8'h9F;
                    16'hA7F9: data_out = 8'hA0;
                    16'hA7FA: data_out = 8'hA1;
                    16'hA7FB: data_out = 8'hA2;
                    16'hA7FC: data_out = 8'hA3;
                    16'hA7FD: data_out = 8'hA4;
                    16'hA7FE: data_out = 8'hA5;
                    16'hA7FF: data_out = 8'hA6;
                    16'hA800: data_out = 8'hA8;
                    16'hA801: data_out = 8'hA7;
                    16'hA802: data_out = 8'hA6;
                    16'hA803: data_out = 8'hA5;
                    16'hA804: data_out = 8'hA4;
                    16'hA805: data_out = 8'hA3;
                    16'hA806: data_out = 8'hA2;
                    16'hA807: data_out = 8'hA1;
                    16'hA808: data_out = 8'hA0;
                    16'hA809: data_out = 8'h9F;
                    16'hA80A: data_out = 8'h9E;
                    16'hA80B: data_out = 8'h9D;
                    16'hA80C: data_out = 8'h9C;
                    16'hA80D: data_out = 8'h9B;
                    16'hA80E: data_out = 8'h9A;
                    16'hA80F: data_out = 8'h99;
                    16'hA810: data_out = 8'h98;
                    16'hA811: data_out = 8'h97;
                    16'hA812: data_out = 8'h96;
                    16'hA813: data_out = 8'h95;
                    16'hA814: data_out = 8'h94;
                    16'hA815: data_out = 8'h93;
                    16'hA816: data_out = 8'h92;
                    16'hA817: data_out = 8'h91;
                    16'hA818: data_out = 8'h90;
                    16'hA819: data_out = 8'h8F;
                    16'hA81A: data_out = 8'h8E;
                    16'hA81B: data_out = 8'h8D;
                    16'hA81C: data_out = 8'h8C;
                    16'hA81D: data_out = 8'h8B;
                    16'hA81E: data_out = 8'h8A;
                    16'hA81F: data_out = 8'h89;
                    16'hA820: data_out = 8'h88;
                    16'hA821: data_out = 8'h87;
                    16'hA822: data_out = 8'h86;
                    16'hA823: data_out = 8'h85;
                    16'hA824: data_out = 8'h84;
                    16'hA825: data_out = 8'h83;
                    16'hA826: data_out = 8'h82;
                    16'hA827: data_out = 8'h81;
                    16'hA828: data_out = 8'h0;
                    16'hA829: data_out = 8'h1;
                    16'hA82A: data_out = 8'h2;
                    16'hA82B: data_out = 8'h3;
                    16'hA82C: data_out = 8'h4;
                    16'hA82D: data_out = 8'h5;
                    16'hA82E: data_out = 8'h6;
                    16'hA82F: data_out = 8'h7;
                    16'hA830: data_out = 8'h8;
                    16'hA831: data_out = 8'h9;
                    16'hA832: data_out = 8'hA;
                    16'hA833: data_out = 8'hB;
                    16'hA834: data_out = 8'hC;
                    16'hA835: data_out = 8'hD;
                    16'hA836: data_out = 8'hE;
                    16'hA837: data_out = 8'hF;
                    16'hA838: data_out = 8'h10;
                    16'hA839: data_out = 8'h11;
                    16'hA83A: data_out = 8'h12;
                    16'hA83B: data_out = 8'h13;
                    16'hA83C: data_out = 8'h14;
                    16'hA83D: data_out = 8'h15;
                    16'hA83E: data_out = 8'h16;
                    16'hA83F: data_out = 8'h17;
                    16'hA840: data_out = 8'h18;
                    16'hA841: data_out = 8'h19;
                    16'hA842: data_out = 8'h1A;
                    16'hA843: data_out = 8'h1B;
                    16'hA844: data_out = 8'h1C;
                    16'hA845: data_out = 8'h1D;
                    16'hA846: data_out = 8'h1E;
                    16'hA847: data_out = 8'h1F;
                    16'hA848: data_out = 8'h20;
                    16'hA849: data_out = 8'h21;
                    16'hA84A: data_out = 8'h22;
                    16'hA84B: data_out = 8'h23;
                    16'hA84C: data_out = 8'h24;
                    16'hA84D: data_out = 8'h25;
                    16'hA84E: data_out = 8'h26;
                    16'hA84F: data_out = 8'h27;
                    16'hA850: data_out = 8'h28;
                    16'hA851: data_out = 8'h29;
                    16'hA852: data_out = 8'h2A;
                    16'hA853: data_out = 8'h2B;
                    16'hA854: data_out = 8'h2C;
                    16'hA855: data_out = 8'h2D;
                    16'hA856: data_out = 8'h2E;
                    16'hA857: data_out = 8'h2F;
                    16'hA858: data_out = 8'h30;
                    16'hA859: data_out = 8'h31;
                    16'hA85A: data_out = 8'h32;
                    16'hA85B: data_out = 8'h33;
                    16'hA85C: data_out = 8'h34;
                    16'hA85D: data_out = 8'h35;
                    16'hA85E: data_out = 8'h36;
                    16'hA85F: data_out = 8'h37;
                    16'hA860: data_out = 8'h38;
                    16'hA861: data_out = 8'h39;
                    16'hA862: data_out = 8'h3A;
                    16'hA863: data_out = 8'h3B;
                    16'hA864: data_out = 8'h3C;
                    16'hA865: data_out = 8'h3D;
                    16'hA866: data_out = 8'h3E;
                    16'hA867: data_out = 8'h3F;
                    16'hA868: data_out = 8'h40;
                    16'hA869: data_out = 8'h41;
                    16'hA86A: data_out = 8'h42;
                    16'hA86B: data_out = 8'h43;
                    16'hA86C: data_out = 8'h44;
                    16'hA86D: data_out = 8'h45;
                    16'hA86E: data_out = 8'h46;
                    16'hA86F: data_out = 8'h47;
                    16'hA870: data_out = 8'h48;
                    16'hA871: data_out = 8'h49;
                    16'hA872: data_out = 8'h4A;
                    16'hA873: data_out = 8'h4B;
                    16'hA874: data_out = 8'h4C;
                    16'hA875: data_out = 8'h4D;
                    16'hA876: data_out = 8'h4E;
                    16'hA877: data_out = 8'h4F;
                    16'hA878: data_out = 8'h50;
                    16'hA879: data_out = 8'h51;
                    16'hA87A: data_out = 8'h52;
                    16'hA87B: data_out = 8'h53;
                    16'hA87C: data_out = 8'h54;
                    16'hA87D: data_out = 8'h55;
                    16'hA87E: data_out = 8'h56;
                    16'hA87F: data_out = 8'h57;
                    16'hA880: data_out = 8'hA8;
                    16'hA881: data_out = 8'hA9;
                    16'hA882: data_out = 8'hAA;
                    16'hA883: data_out = 8'hAB;
                    16'hA884: data_out = 8'hAC;
                    16'hA885: data_out = 8'hAD;
                    16'hA886: data_out = 8'hAE;
                    16'hA887: data_out = 8'hAF;
                    16'hA888: data_out = 8'hB0;
                    16'hA889: data_out = 8'hB1;
                    16'hA88A: data_out = 8'hB2;
                    16'hA88B: data_out = 8'hB3;
                    16'hA88C: data_out = 8'hB4;
                    16'hA88D: data_out = 8'hB5;
                    16'hA88E: data_out = 8'hB6;
                    16'hA88F: data_out = 8'hB7;
                    16'hA890: data_out = 8'hB8;
                    16'hA891: data_out = 8'hB9;
                    16'hA892: data_out = 8'hBA;
                    16'hA893: data_out = 8'hBB;
                    16'hA894: data_out = 8'hBC;
                    16'hA895: data_out = 8'hBD;
                    16'hA896: data_out = 8'hBE;
                    16'hA897: data_out = 8'hBF;
                    16'hA898: data_out = 8'hC0;
                    16'hA899: data_out = 8'hC1;
                    16'hA89A: data_out = 8'hC2;
                    16'hA89B: data_out = 8'hC3;
                    16'hA89C: data_out = 8'hC4;
                    16'hA89D: data_out = 8'hC5;
                    16'hA89E: data_out = 8'hC6;
                    16'hA89F: data_out = 8'hC7;
                    16'hA8A0: data_out = 8'hC8;
                    16'hA8A1: data_out = 8'hC9;
                    16'hA8A2: data_out = 8'hCA;
                    16'hA8A3: data_out = 8'hCB;
                    16'hA8A4: data_out = 8'hCC;
                    16'hA8A5: data_out = 8'hCD;
                    16'hA8A6: data_out = 8'hCE;
                    16'hA8A7: data_out = 8'hCF;
                    16'hA8A8: data_out = 8'hD0;
                    16'hA8A9: data_out = 8'hD1;
                    16'hA8AA: data_out = 8'hD2;
                    16'hA8AB: data_out = 8'hD3;
                    16'hA8AC: data_out = 8'hD4;
                    16'hA8AD: data_out = 8'hD5;
                    16'hA8AE: data_out = 8'hD6;
                    16'hA8AF: data_out = 8'hD7;
                    16'hA8B0: data_out = 8'hD8;
                    16'hA8B1: data_out = 8'hD9;
                    16'hA8B2: data_out = 8'hDA;
                    16'hA8B3: data_out = 8'hDB;
                    16'hA8B4: data_out = 8'hDC;
                    16'hA8B5: data_out = 8'hDD;
                    16'hA8B6: data_out = 8'hDE;
                    16'hA8B7: data_out = 8'hDF;
                    16'hA8B8: data_out = 8'hE0;
                    16'hA8B9: data_out = 8'hE1;
                    16'hA8BA: data_out = 8'hE2;
                    16'hA8BB: data_out = 8'hE3;
                    16'hA8BC: data_out = 8'hE4;
                    16'hA8BD: data_out = 8'hE5;
                    16'hA8BE: data_out = 8'hE6;
                    16'hA8BF: data_out = 8'hE7;
                    16'hA8C0: data_out = 8'hE8;
                    16'hA8C1: data_out = 8'hE9;
                    16'hA8C2: data_out = 8'hEA;
                    16'hA8C3: data_out = 8'hEB;
                    16'hA8C4: data_out = 8'hEC;
                    16'hA8C5: data_out = 8'hED;
                    16'hA8C6: data_out = 8'hEE;
                    16'hA8C7: data_out = 8'hEF;
                    16'hA8C8: data_out = 8'hF0;
                    16'hA8C9: data_out = 8'hF1;
                    16'hA8CA: data_out = 8'hF2;
                    16'hA8CB: data_out = 8'hF3;
                    16'hA8CC: data_out = 8'hF4;
                    16'hA8CD: data_out = 8'hF5;
                    16'hA8CE: data_out = 8'hF6;
                    16'hA8CF: data_out = 8'hF7;
                    16'hA8D0: data_out = 8'hF8;
                    16'hA8D1: data_out = 8'hF9;
                    16'hA8D2: data_out = 8'hFA;
                    16'hA8D3: data_out = 8'hFB;
                    16'hA8D4: data_out = 8'hFC;
                    16'hA8D5: data_out = 8'hFD;
                    16'hA8D6: data_out = 8'hFE;
                    16'hA8D7: data_out = 8'hFF;
                    16'hA8D8: data_out = 8'h80;
                    16'hA8D9: data_out = 8'h81;
                    16'hA8DA: data_out = 8'h82;
                    16'hA8DB: data_out = 8'h83;
                    16'hA8DC: data_out = 8'h84;
                    16'hA8DD: data_out = 8'h85;
                    16'hA8DE: data_out = 8'h86;
                    16'hA8DF: data_out = 8'h87;
                    16'hA8E0: data_out = 8'h88;
                    16'hA8E1: data_out = 8'h89;
                    16'hA8E2: data_out = 8'h8A;
                    16'hA8E3: data_out = 8'h8B;
                    16'hA8E4: data_out = 8'h8C;
                    16'hA8E5: data_out = 8'h8D;
                    16'hA8E6: data_out = 8'h8E;
                    16'hA8E7: data_out = 8'h8F;
                    16'hA8E8: data_out = 8'h90;
                    16'hA8E9: data_out = 8'h91;
                    16'hA8EA: data_out = 8'h92;
                    16'hA8EB: data_out = 8'h93;
                    16'hA8EC: data_out = 8'h94;
                    16'hA8ED: data_out = 8'h95;
                    16'hA8EE: data_out = 8'h96;
                    16'hA8EF: data_out = 8'h97;
                    16'hA8F0: data_out = 8'h98;
                    16'hA8F1: data_out = 8'h99;
                    16'hA8F2: data_out = 8'h9A;
                    16'hA8F3: data_out = 8'h9B;
                    16'hA8F4: data_out = 8'h9C;
                    16'hA8F5: data_out = 8'h9D;
                    16'hA8F6: data_out = 8'h9E;
                    16'hA8F7: data_out = 8'h9F;
                    16'hA8F8: data_out = 8'hA0;
                    16'hA8F9: data_out = 8'hA1;
                    16'hA8FA: data_out = 8'hA2;
                    16'hA8FB: data_out = 8'hA3;
                    16'hA8FC: data_out = 8'hA4;
                    16'hA8FD: data_out = 8'hA5;
                    16'hA8FE: data_out = 8'hA6;
                    16'hA8FF: data_out = 8'hA7;
                    16'hA900: data_out = 8'hA9;
                    16'hA901: data_out = 8'hA8;
                    16'hA902: data_out = 8'hA7;
                    16'hA903: data_out = 8'hA6;
                    16'hA904: data_out = 8'hA5;
                    16'hA905: data_out = 8'hA4;
                    16'hA906: data_out = 8'hA3;
                    16'hA907: data_out = 8'hA2;
                    16'hA908: data_out = 8'hA1;
                    16'hA909: data_out = 8'hA0;
                    16'hA90A: data_out = 8'h9F;
                    16'hA90B: data_out = 8'h9E;
                    16'hA90C: data_out = 8'h9D;
                    16'hA90D: data_out = 8'h9C;
                    16'hA90E: data_out = 8'h9B;
                    16'hA90F: data_out = 8'h9A;
                    16'hA910: data_out = 8'h99;
                    16'hA911: data_out = 8'h98;
                    16'hA912: data_out = 8'h97;
                    16'hA913: data_out = 8'h96;
                    16'hA914: data_out = 8'h95;
                    16'hA915: data_out = 8'h94;
                    16'hA916: data_out = 8'h93;
                    16'hA917: data_out = 8'h92;
                    16'hA918: data_out = 8'h91;
                    16'hA919: data_out = 8'h90;
                    16'hA91A: data_out = 8'h8F;
                    16'hA91B: data_out = 8'h8E;
                    16'hA91C: data_out = 8'h8D;
                    16'hA91D: data_out = 8'h8C;
                    16'hA91E: data_out = 8'h8B;
                    16'hA91F: data_out = 8'h8A;
                    16'hA920: data_out = 8'h89;
                    16'hA921: data_out = 8'h88;
                    16'hA922: data_out = 8'h87;
                    16'hA923: data_out = 8'h86;
                    16'hA924: data_out = 8'h85;
                    16'hA925: data_out = 8'h84;
                    16'hA926: data_out = 8'h83;
                    16'hA927: data_out = 8'h82;
                    16'hA928: data_out = 8'h81;
                    16'hA929: data_out = 8'h0;
                    16'hA92A: data_out = 8'h1;
                    16'hA92B: data_out = 8'h2;
                    16'hA92C: data_out = 8'h3;
                    16'hA92D: data_out = 8'h4;
                    16'hA92E: data_out = 8'h5;
                    16'hA92F: data_out = 8'h6;
                    16'hA930: data_out = 8'h7;
                    16'hA931: data_out = 8'h8;
                    16'hA932: data_out = 8'h9;
                    16'hA933: data_out = 8'hA;
                    16'hA934: data_out = 8'hB;
                    16'hA935: data_out = 8'hC;
                    16'hA936: data_out = 8'hD;
                    16'hA937: data_out = 8'hE;
                    16'hA938: data_out = 8'hF;
                    16'hA939: data_out = 8'h10;
                    16'hA93A: data_out = 8'h11;
                    16'hA93B: data_out = 8'h12;
                    16'hA93C: data_out = 8'h13;
                    16'hA93D: data_out = 8'h14;
                    16'hA93E: data_out = 8'h15;
                    16'hA93F: data_out = 8'h16;
                    16'hA940: data_out = 8'h17;
                    16'hA941: data_out = 8'h18;
                    16'hA942: data_out = 8'h19;
                    16'hA943: data_out = 8'h1A;
                    16'hA944: data_out = 8'h1B;
                    16'hA945: data_out = 8'h1C;
                    16'hA946: data_out = 8'h1D;
                    16'hA947: data_out = 8'h1E;
                    16'hA948: data_out = 8'h1F;
                    16'hA949: data_out = 8'h20;
                    16'hA94A: data_out = 8'h21;
                    16'hA94B: data_out = 8'h22;
                    16'hA94C: data_out = 8'h23;
                    16'hA94D: data_out = 8'h24;
                    16'hA94E: data_out = 8'h25;
                    16'hA94F: data_out = 8'h26;
                    16'hA950: data_out = 8'h27;
                    16'hA951: data_out = 8'h28;
                    16'hA952: data_out = 8'h29;
                    16'hA953: data_out = 8'h2A;
                    16'hA954: data_out = 8'h2B;
                    16'hA955: data_out = 8'h2C;
                    16'hA956: data_out = 8'h2D;
                    16'hA957: data_out = 8'h2E;
                    16'hA958: data_out = 8'h2F;
                    16'hA959: data_out = 8'h30;
                    16'hA95A: data_out = 8'h31;
                    16'hA95B: data_out = 8'h32;
                    16'hA95C: data_out = 8'h33;
                    16'hA95D: data_out = 8'h34;
                    16'hA95E: data_out = 8'h35;
                    16'hA95F: data_out = 8'h36;
                    16'hA960: data_out = 8'h37;
                    16'hA961: data_out = 8'h38;
                    16'hA962: data_out = 8'h39;
                    16'hA963: data_out = 8'h3A;
                    16'hA964: data_out = 8'h3B;
                    16'hA965: data_out = 8'h3C;
                    16'hA966: data_out = 8'h3D;
                    16'hA967: data_out = 8'h3E;
                    16'hA968: data_out = 8'h3F;
                    16'hA969: data_out = 8'h40;
                    16'hA96A: data_out = 8'h41;
                    16'hA96B: data_out = 8'h42;
                    16'hA96C: data_out = 8'h43;
                    16'hA96D: data_out = 8'h44;
                    16'hA96E: data_out = 8'h45;
                    16'hA96F: data_out = 8'h46;
                    16'hA970: data_out = 8'h47;
                    16'hA971: data_out = 8'h48;
                    16'hA972: data_out = 8'h49;
                    16'hA973: data_out = 8'h4A;
                    16'hA974: data_out = 8'h4B;
                    16'hA975: data_out = 8'h4C;
                    16'hA976: data_out = 8'h4D;
                    16'hA977: data_out = 8'h4E;
                    16'hA978: data_out = 8'h4F;
                    16'hA979: data_out = 8'h50;
                    16'hA97A: data_out = 8'h51;
                    16'hA97B: data_out = 8'h52;
                    16'hA97C: data_out = 8'h53;
                    16'hA97D: data_out = 8'h54;
                    16'hA97E: data_out = 8'h55;
                    16'hA97F: data_out = 8'h56;
                    16'hA980: data_out = 8'hA9;
                    16'hA981: data_out = 8'hAA;
                    16'hA982: data_out = 8'hAB;
                    16'hA983: data_out = 8'hAC;
                    16'hA984: data_out = 8'hAD;
                    16'hA985: data_out = 8'hAE;
                    16'hA986: data_out = 8'hAF;
                    16'hA987: data_out = 8'hB0;
                    16'hA988: data_out = 8'hB1;
                    16'hA989: data_out = 8'hB2;
                    16'hA98A: data_out = 8'hB3;
                    16'hA98B: data_out = 8'hB4;
                    16'hA98C: data_out = 8'hB5;
                    16'hA98D: data_out = 8'hB6;
                    16'hA98E: data_out = 8'hB7;
                    16'hA98F: data_out = 8'hB8;
                    16'hA990: data_out = 8'hB9;
                    16'hA991: data_out = 8'hBA;
                    16'hA992: data_out = 8'hBB;
                    16'hA993: data_out = 8'hBC;
                    16'hA994: data_out = 8'hBD;
                    16'hA995: data_out = 8'hBE;
                    16'hA996: data_out = 8'hBF;
                    16'hA997: data_out = 8'hC0;
                    16'hA998: data_out = 8'hC1;
                    16'hA999: data_out = 8'hC2;
                    16'hA99A: data_out = 8'hC3;
                    16'hA99B: data_out = 8'hC4;
                    16'hA99C: data_out = 8'hC5;
                    16'hA99D: data_out = 8'hC6;
                    16'hA99E: data_out = 8'hC7;
                    16'hA99F: data_out = 8'hC8;
                    16'hA9A0: data_out = 8'hC9;
                    16'hA9A1: data_out = 8'hCA;
                    16'hA9A2: data_out = 8'hCB;
                    16'hA9A3: data_out = 8'hCC;
                    16'hA9A4: data_out = 8'hCD;
                    16'hA9A5: data_out = 8'hCE;
                    16'hA9A6: data_out = 8'hCF;
                    16'hA9A7: data_out = 8'hD0;
                    16'hA9A8: data_out = 8'hD1;
                    16'hA9A9: data_out = 8'hD2;
                    16'hA9AA: data_out = 8'hD3;
                    16'hA9AB: data_out = 8'hD4;
                    16'hA9AC: data_out = 8'hD5;
                    16'hA9AD: data_out = 8'hD6;
                    16'hA9AE: data_out = 8'hD7;
                    16'hA9AF: data_out = 8'hD8;
                    16'hA9B0: data_out = 8'hD9;
                    16'hA9B1: data_out = 8'hDA;
                    16'hA9B2: data_out = 8'hDB;
                    16'hA9B3: data_out = 8'hDC;
                    16'hA9B4: data_out = 8'hDD;
                    16'hA9B5: data_out = 8'hDE;
                    16'hA9B6: data_out = 8'hDF;
                    16'hA9B7: data_out = 8'hE0;
                    16'hA9B8: data_out = 8'hE1;
                    16'hA9B9: data_out = 8'hE2;
                    16'hA9BA: data_out = 8'hE3;
                    16'hA9BB: data_out = 8'hE4;
                    16'hA9BC: data_out = 8'hE5;
                    16'hA9BD: data_out = 8'hE6;
                    16'hA9BE: data_out = 8'hE7;
                    16'hA9BF: data_out = 8'hE8;
                    16'hA9C0: data_out = 8'hE9;
                    16'hA9C1: data_out = 8'hEA;
                    16'hA9C2: data_out = 8'hEB;
                    16'hA9C3: data_out = 8'hEC;
                    16'hA9C4: data_out = 8'hED;
                    16'hA9C5: data_out = 8'hEE;
                    16'hA9C6: data_out = 8'hEF;
                    16'hA9C7: data_out = 8'hF0;
                    16'hA9C8: data_out = 8'hF1;
                    16'hA9C9: data_out = 8'hF2;
                    16'hA9CA: data_out = 8'hF3;
                    16'hA9CB: data_out = 8'hF4;
                    16'hA9CC: data_out = 8'hF5;
                    16'hA9CD: data_out = 8'hF6;
                    16'hA9CE: data_out = 8'hF7;
                    16'hA9CF: data_out = 8'hF8;
                    16'hA9D0: data_out = 8'hF9;
                    16'hA9D1: data_out = 8'hFA;
                    16'hA9D2: data_out = 8'hFB;
                    16'hA9D3: data_out = 8'hFC;
                    16'hA9D4: data_out = 8'hFD;
                    16'hA9D5: data_out = 8'hFE;
                    16'hA9D6: data_out = 8'hFF;
                    16'hA9D7: data_out = 8'h80;
                    16'hA9D8: data_out = 8'h81;
                    16'hA9D9: data_out = 8'h82;
                    16'hA9DA: data_out = 8'h83;
                    16'hA9DB: data_out = 8'h84;
                    16'hA9DC: data_out = 8'h85;
                    16'hA9DD: data_out = 8'h86;
                    16'hA9DE: data_out = 8'h87;
                    16'hA9DF: data_out = 8'h88;
                    16'hA9E0: data_out = 8'h89;
                    16'hA9E1: data_out = 8'h8A;
                    16'hA9E2: data_out = 8'h8B;
                    16'hA9E3: data_out = 8'h8C;
                    16'hA9E4: data_out = 8'h8D;
                    16'hA9E5: data_out = 8'h8E;
                    16'hA9E6: data_out = 8'h8F;
                    16'hA9E7: data_out = 8'h90;
                    16'hA9E8: data_out = 8'h91;
                    16'hA9E9: data_out = 8'h92;
                    16'hA9EA: data_out = 8'h93;
                    16'hA9EB: data_out = 8'h94;
                    16'hA9EC: data_out = 8'h95;
                    16'hA9ED: data_out = 8'h96;
                    16'hA9EE: data_out = 8'h97;
                    16'hA9EF: data_out = 8'h98;
                    16'hA9F0: data_out = 8'h99;
                    16'hA9F1: data_out = 8'h9A;
                    16'hA9F2: data_out = 8'h9B;
                    16'hA9F3: data_out = 8'h9C;
                    16'hA9F4: data_out = 8'h9D;
                    16'hA9F5: data_out = 8'h9E;
                    16'hA9F6: data_out = 8'h9F;
                    16'hA9F7: data_out = 8'hA0;
                    16'hA9F8: data_out = 8'hA1;
                    16'hA9F9: data_out = 8'hA2;
                    16'hA9FA: data_out = 8'hA3;
                    16'hA9FB: data_out = 8'hA4;
                    16'hA9FC: data_out = 8'hA5;
                    16'hA9FD: data_out = 8'hA6;
                    16'hA9FE: data_out = 8'hA7;
                    16'hA9FF: data_out = 8'hA8;
                    16'hAA00: data_out = 8'hAA;
                    16'hAA01: data_out = 8'hA9;
                    16'hAA02: data_out = 8'hA8;
                    16'hAA03: data_out = 8'hA7;
                    16'hAA04: data_out = 8'hA6;
                    16'hAA05: data_out = 8'hA5;
                    16'hAA06: data_out = 8'hA4;
                    16'hAA07: data_out = 8'hA3;
                    16'hAA08: data_out = 8'hA2;
                    16'hAA09: data_out = 8'hA1;
                    16'hAA0A: data_out = 8'hA0;
                    16'hAA0B: data_out = 8'h9F;
                    16'hAA0C: data_out = 8'h9E;
                    16'hAA0D: data_out = 8'h9D;
                    16'hAA0E: data_out = 8'h9C;
                    16'hAA0F: data_out = 8'h9B;
                    16'hAA10: data_out = 8'h9A;
                    16'hAA11: data_out = 8'h99;
                    16'hAA12: data_out = 8'h98;
                    16'hAA13: data_out = 8'h97;
                    16'hAA14: data_out = 8'h96;
                    16'hAA15: data_out = 8'h95;
                    16'hAA16: data_out = 8'h94;
                    16'hAA17: data_out = 8'h93;
                    16'hAA18: data_out = 8'h92;
                    16'hAA19: data_out = 8'h91;
                    16'hAA1A: data_out = 8'h90;
                    16'hAA1B: data_out = 8'h8F;
                    16'hAA1C: data_out = 8'h8E;
                    16'hAA1D: data_out = 8'h8D;
                    16'hAA1E: data_out = 8'h8C;
                    16'hAA1F: data_out = 8'h8B;
                    16'hAA20: data_out = 8'h8A;
                    16'hAA21: data_out = 8'h89;
                    16'hAA22: data_out = 8'h88;
                    16'hAA23: data_out = 8'h87;
                    16'hAA24: data_out = 8'h86;
                    16'hAA25: data_out = 8'h85;
                    16'hAA26: data_out = 8'h84;
                    16'hAA27: data_out = 8'h83;
                    16'hAA28: data_out = 8'h82;
                    16'hAA29: data_out = 8'h81;
                    16'hAA2A: data_out = 8'h0;
                    16'hAA2B: data_out = 8'h1;
                    16'hAA2C: data_out = 8'h2;
                    16'hAA2D: data_out = 8'h3;
                    16'hAA2E: data_out = 8'h4;
                    16'hAA2F: data_out = 8'h5;
                    16'hAA30: data_out = 8'h6;
                    16'hAA31: data_out = 8'h7;
                    16'hAA32: data_out = 8'h8;
                    16'hAA33: data_out = 8'h9;
                    16'hAA34: data_out = 8'hA;
                    16'hAA35: data_out = 8'hB;
                    16'hAA36: data_out = 8'hC;
                    16'hAA37: data_out = 8'hD;
                    16'hAA38: data_out = 8'hE;
                    16'hAA39: data_out = 8'hF;
                    16'hAA3A: data_out = 8'h10;
                    16'hAA3B: data_out = 8'h11;
                    16'hAA3C: data_out = 8'h12;
                    16'hAA3D: data_out = 8'h13;
                    16'hAA3E: data_out = 8'h14;
                    16'hAA3F: data_out = 8'h15;
                    16'hAA40: data_out = 8'h16;
                    16'hAA41: data_out = 8'h17;
                    16'hAA42: data_out = 8'h18;
                    16'hAA43: data_out = 8'h19;
                    16'hAA44: data_out = 8'h1A;
                    16'hAA45: data_out = 8'h1B;
                    16'hAA46: data_out = 8'h1C;
                    16'hAA47: data_out = 8'h1D;
                    16'hAA48: data_out = 8'h1E;
                    16'hAA49: data_out = 8'h1F;
                    16'hAA4A: data_out = 8'h20;
                    16'hAA4B: data_out = 8'h21;
                    16'hAA4C: data_out = 8'h22;
                    16'hAA4D: data_out = 8'h23;
                    16'hAA4E: data_out = 8'h24;
                    16'hAA4F: data_out = 8'h25;
                    16'hAA50: data_out = 8'h26;
                    16'hAA51: data_out = 8'h27;
                    16'hAA52: data_out = 8'h28;
                    16'hAA53: data_out = 8'h29;
                    16'hAA54: data_out = 8'h2A;
                    16'hAA55: data_out = 8'h2B;
                    16'hAA56: data_out = 8'h2C;
                    16'hAA57: data_out = 8'h2D;
                    16'hAA58: data_out = 8'h2E;
                    16'hAA59: data_out = 8'h2F;
                    16'hAA5A: data_out = 8'h30;
                    16'hAA5B: data_out = 8'h31;
                    16'hAA5C: data_out = 8'h32;
                    16'hAA5D: data_out = 8'h33;
                    16'hAA5E: data_out = 8'h34;
                    16'hAA5F: data_out = 8'h35;
                    16'hAA60: data_out = 8'h36;
                    16'hAA61: data_out = 8'h37;
                    16'hAA62: data_out = 8'h38;
                    16'hAA63: data_out = 8'h39;
                    16'hAA64: data_out = 8'h3A;
                    16'hAA65: data_out = 8'h3B;
                    16'hAA66: data_out = 8'h3C;
                    16'hAA67: data_out = 8'h3D;
                    16'hAA68: data_out = 8'h3E;
                    16'hAA69: data_out = 8'h3F;
                    16'hAA6A: data_out = 8'h40;
                    16'hAA6B: data_out = 8'h41;
                    16'hAA6C: data_out = 8'h42;
                    16'hAA6D: data_out = 8'h43;
                    16'hAA6E: data_out = 8'h44;
                    16'hAA6F: data_out = 8'h45;
                    16'hAA70: data_out = 8'h46;
                    16'hAA71: data_out = 8'h47;
                    16'hAA72: data_out = 8'h48;
                    16'hAA73: data_out = 8'h49;
                    16'hAA74: data_out = 8'h4A;
                    16'hAA75: data_out = 8'h4B;
                    16'hAA76: data_out = 8'h4C;
                    16'hAA77: data_out = 8'h4D;
                    16'hAA78: data_out = 8'h4E;
                    16'hAA79: data_out = 8'h4F;
                    16'hAA7A: data_out = 8'h50;
                    16'hAA7B: data_out = 8'h51;
                    16'hAA7C: data_out = 8'h52;
                    16'hAA7D: data_out = 8'h53;
                    16'hAA7E: data_out = 8'h54;
                    16'hAA7F: data_out = 8'h55;
                    16'hAA80: data_out = 8'hAA;
                    16'hAA81: data_out = 8'hAB;
                    16'hAA82: data_out = 8'hAC;
                    16'hAA83: data_out = 8'hAD;
                    16'hAA84: data_out = 8'hAE;
                    16'hAA85: data_out = 8'hAF;
                    16'hAA86: data_out = 8'hB0;
                    16'hAA87: data_out = 8'hB1;
                    16'hAA88: data_out = 8'hB2;
                    16'hAA89: data_out = 8'hB3;
                    16'hAA8A: data_out = 8'hB4;
                    16'hAA8B: data_out = 8'hB5;
                    16'hAA8C: data_out = 8'hB6;
                    16'hAA8D: data_out = 8'hB7;
                    16'hAA8E: data_out = 8'hB8;
                    16'hAA8F: data_out = 8'hB9;
                    16'hAA90: data_out = 8'hBA;
                    16'hAA91: data_out = 8'hBB;
                    16'hAA92: data_out = 8'hBC;
                    16'hAA93: data_out = 8'hBD;
                    16'hAA94: data_out = 8'hBE;
                    16'hAA95: data_out = 8'hBF;
                    16'hAA96: data_out = 8'hC0;
                    16'hAA97: data_out = 8'hC1;
                    16'hAA98: data_out = 8'hC2;
                    16'hAA99: data_out = 8'hC3;
                    16'hAA9A: data_out = 8'hC4;
                    16'hAA9B: data_out = 8'hC5;
                    16'hAA9C: data_out = 8'hC6;
                    16'hAA9D: data_out = 8'hC7;
                    16'hAA9E: data_out = 8'hC8;
                    16'hAA9F: data_out = 8'hC9;
                    16'hAAA0: data_out = 8'hCA;
                    16'hAAA1: data_out = 8'hCB;
                    16'hAAA2: data_out = 8'hCC;
                    16'hAAA3: data_out = 8'hCD;
                    16'hAAA4: data_out = 8'hCE;
                    16'hAAA5: data_out = 8'hCF;
                    16'hAAA6: data_out = 8'hD0;
                    16'hAAA7: data_out = 8'hD1;
                    16'hAAA8: data_out = 8'hD2;
                    16'hAAA9: data_out = 8'hD3;
                    16'hAAAA: data_out = 8'hD4;
                    16'hAAAB: data_out = 8'hD5;
                    16'hAAAC: data_out = 8'hD6;
                    16'hAAAD: data_out = 8'hD7;
                    16'hAAAE: data_out = 8'hD8;
                    16'hAAAF: data_out = 8'hD9;
                    16'hAAB0: data_out = 8'hDA;
                    16'hAAB1: data_out = 8'hDB;
                    16'hAAB2: data_out = 8'hDC;
                    16'hAAB3: data_out = 8'hDD;
                    16'hAAB4: data_out = 8'hDE;
                    16'hAAB5: data_out = 8'hDF;
                    16'hAAB6: data_out = 8'hE0;
                    16'hAAB7: data_out = 8'hE1;
                    16'hAAB8: data_out = 8'hE2;
                    16'hAAB9: data_out = 8'hE3;
                    16'hAABA: data_out = 8'hE4;
                    16'hAABB: data_out = 8'hE5;
                    16'hAABC: data_out = 8'hE6;
                    16'hAABD: data_out = 8'hE7;
                    16'hAABE: data_out = 8'hE8;
                    16'hAABF: data_out = 8'hE9;
                    16'hAAC0: data_out = 8'hEA;
                    16'hAAC1: data_out = 8'hEB;
                    16'hAAC2: data_out = 8'hEC;
                    16'hAAC3: data_out = 8'hED;
                    16'hAAC4: data_out = 8'hEE;
                    16'hAAC5: data_out = 8'hEF;
                    16'hAAC6: data_out = 8'hF0;
                    16'hAAC7: data_out = 8'hF1;
                    16'hAAC8: data_out = 8'hF2;
                    16'hAAC9: data_out = 8'hF3;
                    16'hAACA: data_out = 8'hF4;
                    16'hAACB: data_out = 8'hF5;
                    16'hAACC: data_out = 8'hF6;
                    16'hAACD: data_out = 8'hF7;
                    16'hAACE: data_out = 8'hF8;
                    16'hAACF: data_out = 8'hF9;
                    16'hAAD0: data_out = 8'hFA;
                    16'hAAD1: data_out = 8'hFB;
                    16'hAAD2: data_out = 8'hFC;
                    16'hAAD3: data_out = 8'hFD;
                    16'hAAD4: data_out = 8'hFE;
                    16'hAAD5: data_out = 8'hFF;
                    16'hAAD6: data_out = 8'h80;
                    16'hAAD7: data_out = 8'h81;
                    16'hAAD8: data_out = 8'h82;
                    16'hAAD9: data_out = 8'h83;
                    16'hAADA: data_out = 8'h84;
                    16'hAADB: data_out = 8'h85;
                    16'hAADC: data_out = 8'h86;
                    16'hAADD: data_out = 8'h87;
                    16'hAADE: data_out = 8'h88;
                    16'hAADF: data_out = 8'h89;
                    16'hAAE0: data_out = 8'h8A;
                    16'hAAE1: data_out = 8'h8B;
                    16'hAAE2: data_out = 8'h8C;
                    16'hAAE3: data_out = 8'h8D;
                    16'hAAE4: data_out = 8'h8E;
                    16'hAAE5: data_out = 8'h8F;
                    16'hAAE6: data_out = 8'h90;
                    16'hAAE7: data_out = 8'h91;
                    16'hAAE8: data_out = 8'h92;
                    16'hAAE9: data_out = 8'h93;
                    16'hAAEA: data_out = 8'h94;
                    16'hAAEB: data_out = 8'h95;
                    16'hAAEC: data_out = 8'h96;
                    16'hAAED: data_out = 8'h97;
                    16'hAAEE: data_out = 8'h98;
                    16'hAAEF: data_out = 8'h99;
                    16'hAAF0: data_out = 8'h9A;
                    16'hAAF1: data_out = 8'h9B;
                    16'hAAF2: data_out = 8'h9C;
                    16'hAAF3: data_out = 8'h9D;
                    16'hAAF4: data_out = 8'h9E;
                    16'hAAF5: data_out = 8'h9F;
                    16'hAAF6: data_out = 8'hA0;
                    16'hAAF7: data_out = 8'hA1;
                    16'hAAF8: data_out = 8'hA2;
                    16'hAAF9: data_out = 8'hA3;
                    16'hAAFA: data_out = 8'hA4;
                    16'hAAFB: data_out = 8'hA5;
                    16'hAAFC: data_out = 8'hA6;
                    16'hAAFD: data_out = 8'hA7;
                    16'hAAFE: data_out = 8'hA8;
                    16'hAAFF: data_out = 8'hA9;
                    16'hAB00: data_out = 8'hAB;
                    16'hAB01: data_out = 8'hAA;
                    16'hAB02: data_out = 8'hA9;
                    16'hAB03: data_out = 8'hA8;
                    16'hAB04: data_out = 8'hA7;
                    16'hAB05: data_out = 8'hA6;
                    16'hAB06: data_out = 8'hA5;
                    16'hAB07: data_out = 8'hA4;
                    16'hAB08: data_out = 8'hA3;
                    16'hAB09: data_out = 8'hA2;
                    16'hAB0A: data_out = 8'hA1;
                    16'hAB0B: data_out = 8'hA0;
                    16'hAB0C: data_out = 8'h9F;
                    16'hAB0D: data_out = 8'h9E;
                    16'hAB0E: data_out = 8'h9D;
                    16'hAB0F: data_out = 8'h9C;
                    16'hAB10: data_out = 8'h9B;
                    16'hAB11: data_out = 8'h9A;
                    16'hAB12: data_out = 8'h99;
                    16'hAB13: data_out = 8'h98;
                    16'hAB14: data_out = 8'h97;
                    16'hAB15: data_out = 8'h96;
                    16'hAB16: data_out = 8'h95;
                    16'hAB17: data_out = 8'h94;
                    16'hAB18: data_out = 8'h93;
                    16'hAB19: data_out = 8'h92;
                    16'hAB1A: data_out = 8'h91;
                    16'hAB1B: data_out = 8'h90;
                    16'hAB1C: data_out = 8'h8F;
                    16'hAB1D: data_out = 8'h8E;
                    16'hAB1E: data_out = 8'h8D;
                    16'hAB1F: data_out = 8'h8C;
                    16'hAB20: data_out = 8'h8B;
                    16'hAB21: data_out = 8'h8A;
                    16'hAB22: data_out = 8'h89;
                    16'hAB23: data_out = 8'h88;
                    16'hAB24: data_out = 8'h87;
                    16'hAB25: data_out = 8'h86;
                    16'hAB26: data_out = 8'h85;
                    16'hAB27: data_out = 8'h84;
                    16'hAB28: data_out = 8'h83;
                    16'hAB29: data_out = 8'h82;
                    16'hAB2A: data_out = 8'h81;
                    16'hAB2B: data_out = 8'h0;
                    16'hAB2C: data_out = 8'h1;
                    16'hAB2D: data_out = 8'h2;
                    16'hAB2E: data_out = 8'h3;
                    16'hAB2F: data_out = 8'h4;
                    16'hAB30: data_out = 8'h5;
                    16'hAB31: data_out = 8'h6;
                    16'hAB32: data_out = 8'h7;
                    16'hAB33: data_out = 8'h8;
                    16'hAB34: data_out = 8'h9;
                    16'hAB35: data_out = 8'hA;
                    16'hAB36: data_out = 8'hB;
                    16'hAB37: data_out = 8'hC;
                    16'hAB38: data_out = 8'hD;
                    16'hAB39: data_out = 8'hE;
                    16'hAB3A: data_out = 8'hF;
                    16'hAB3B: data_out = 8'h10;
                    16'hAB3C: data_out = 8'h11;
                    16'hAB3D: data_out = 8'h12;
                    16'hAB3E: data_out = 8'h13;
                    16'hAB3F: data_out = 8'h14;
                    16'hAB40: data_out = 8'h15;
                    16'hAB41: data_out = 8'h16;
                    16'hAB42: data_out = 8'h17;
                    16'hAB43: data_out = 8'h18;
                    16'hAB44: data_out = 8'h19;
                    16'hAB45: data_out = 8'h1A;
                    16'hAB46: data_out = 8'h1B;
                    16'hAB47: data_out = 8'h1C;
                    16'hAB48: data_out = 8'h1D;
                    16'hAB49: data_out = 8'h1E;
                    16'hAB4A: data_out = 8'h1F;
                    16'hAB4B: data_out = 8'h20;
                    16'hAB4C: data_out = 8'h21;
                    16'hAB4D: data_out = 8'h22;
                    16'hAB4E: data_out = 8'h23;
                    16'hAB4F: data_out = 8'h24;
                    16'hAB50: data_out = 8'h25;
                    16'hAB51: data_out = 8'h26;
                    16'hAB52: data_out = 8'h27;
                    16'hAB53: data_out = 8'h28;
                    16'hAB54: data_out = 8'h29;
                    16'hAB55: data_out = 8'h2A;
                    16'hAB56: data_out = 8'h2B;
                    16'hAB57: data_out = 8'h2C;
                    16'hAB58: data_out = 8'h2D;
                    16'hAB59: data_out = 8'h2E;
                    16'hAB5A: data_out = 8'h2F;
                    16'hAB5B: data_out = 8'h30;
                    16'hAB5C: data_out = 8'h31;
                    16'hAB5D: data_out = 8'h32;
                    16'hAB5E: data_out = 8'h33;
                    16'hAB5F: data_out = 8'h34;
                    16'hAB60: data_out = 8'h35;
                    16'hAB61: data_out = 8'h36;
                    16'hAB62: data_out = 8'h37;
                    16'hAB63: data_out = 8'h38;
                    16'hAB64: data_out = 8'h39;
                    16'hAB65: data_out = 8'h3A;
                    16'hAB66: data_out = 8'h3B;
                    16'hAB67: data_out = 8'h3C;
                    16'hAB68: data_out = 8'h3D;
                    16'hAB69: data_out = 8'h3E;
                    16'hAB6A: data_out = 8'h3F;
                    16'hAB6B: data_out = 8'h40;
                    16'hAB6C: data_out = 8'h41;
                    16'hAB6D: data_out = 8'h42;
                    16'hAB6E: data_out = 8'h43;
                    16'hAB6F: data_out = 8'h44;
                    16'hAB70: data_out = 8'h45;
                    16'hAB71: data_out = 8'h46;
                    16'hAB72: data_out = 8'h47;
                    16'hAB73: data_out = 8'h48;
                    16'hAB74: data_out = 8'h49;
                    16'hAB75: data_out = 8'h4A;
                    16'hAB76: data_out = 8'h4B;
                    16'hAB77: data_out = 8'h4C;
                    16'hAB78: data_out = 8'h4D;
                    16'hAB79: data_out = 8'h4E;
                    16'hAB7A: data_out = 8'h4F;
                    16'hAB7B: data_out = 8'h50;
                    16'hAB7C: data_out = 8'h51;
                    16'hAB7D: data_out = 8'h52;
                    16'hAB7E: data_out = 8'h53;
                    16'hAB7F: data_out = 8'h54;
                    16'hAB80: data_out = 8'hAB;
                    16'hAB81: data_out = 8'hAC;
                    16'hAB82: data_out = 8'hAD;
                    16'hAB83: data_out = 8'hAE;
                    16'hAB84: data_out = 8'hAF;
                    16'hAB85: data_out = 8'hB0;
                    16'hAB86: data_out = 8'hB1;
                    16'hAB87: data_out = 8'hB2;
                    16'hAB88: data_out = 8'hB3;
                    16'hAB89: data_out = 8'hB4;
                    16'hAB8A: data_out = 8'hB5;
                    16'hAB8B: data_out = 8'hB6;
                    16'hAB8C: data_out = 8'hB7;
                    16'hAB8D: data_out = 8'hB8;
                    16'hAB8E: data_out = 8'hB9;
                    16'hAB8F: data_out = 8'hBA;
                    16'hAB90: data_out = 8'hBB;
                    16'hAB91: data_out = 8'hBC;
                    16'hAB92: data_out = 8'hBD;
                    16'hAB93: data_out = 8'hBE;
                    16'hAB94: data_out = 8'hBF;
                    16'hAB95: data_out = 8'hC0;
                    16'hAB96: data_out = 8'hC1;
                    16'hAB97: data_out = 8'hC2;
                    16'hAB98: data_out = 8'hC3;
                    16'hAB99: data_out = 8'hC4;
                    16'hAB9A: data_out = 8'hC5;
                    16'hAB9B: data_out = 8'hC6;
                    16'hAB9C: data_out = 8'hC7;
                    16'hAB9D: data_out = 8'hC8;
                    16'hAB9E: data_out = 8'hC9;
                    16'hAB9F: data_out = 8'hCA;
                    16'hABA0: data_out = 8'hCB;
                    16'hABA1: data_out = 8'hCC;
                    16'hABA2: data_out = 8'hCD;
                    16'hABA3: data_out = 8'hCE;
                    16'hABA4: data_out = 8'hCF;
                    16'hABA5: data_out = 8'hD0;
                    16'hABA6: data_out = 8'hD1;
                    16'hABA7: data_out = 8'hD2;
                    16'hABA8: data_out = 8'hD3;
                    16'hABA9: data_out = 8'hD4;
                    16'hABAA: data_out = 8'hD5;
                    16'hABAB: data_out = 8'hD6;
                    16'hABAC: data_out = 8'hD7;
                    16'hABAD: data_out = 8'hD8;
                    16'hABAE: data_out = 8'hD9;
                    16'hABAF: data_out = 8'hDA;
                    16'hABB0: data_out = 8'hDB;
                    16'hABB1: data_out = 8'hDC;
                    16'hABB2: data_out = 8'hDD;
                    16'hABB3: data_out = 8'hDE;
                    16'hABB4: data_out = 8'hDF;
                    16'hABB5: data_out = 8'hE0;
                    16'hABB6: data_out = 8'hE1;
                    16'hABB7: data_out = 8'hE2;
                    16'hABB8: data_out = 8'hE3;
                    16'hABB9: data_out = 8'hE4;
                    16'hABBA: data_out = 8'hE5;
                    16'hABBB: data_out = 8'hE6;
                    16'hABBC: data_out = 8'hE7;
                    16'hABBD: data_out = 8'hE8;
                    16'hABBE: data_out = 8'hE9;
                    16'hABBF: data_out = 8'hEA;
                    16'hABC0: data_out = 8'hEB;
                    16'hABC1: data_out = 8'hEC;
                    16'hABC2: data_out = 8'hED;
                    16'hABC3: data_out = 8'hEE;
                    16'hABC4: data_out = 8'hEF;
                    16'hABC5: data_out = 8'hF0;
                    16'hABC6: data_out = 8'hF1;
                    16'hABC7: data_out = 8'hF2;
                    16'hABC8: data_out = 8'hF3;
                    16'hABC9: data_out = 8'hF4;
                    16'hABCA: data_out = 8'hF5;
                    16'hABCB: data_out = 8'hF6;
                    16'hABCC: data_out = 8'hF7;
                    16'hABCD: data_out = 8'hF8;
                    16'hABCE: data_out = 8'hF9;
                    16'hABCF: data_out = 8'hFA;
                    16'hABD0: data_out = 8'hFB;
                    16'hABD1: data_out = 8'hFC;
                    16'hABD2: data_out = 8'hFD;
                    16'hABD3: data_out = 8'hFE;
                    16'hABD4: data_out = 8'hFF;
                    16'hABD5: data_out = 8'h80;
                    16'hABD6: data_out = 8'h81;
                    16'hABD7: data_out = 8'h82;
                    16'hABD8: data_out = 8'h83;
                    16'hABD9: data_out = 8'h84;
                    16'hABDA: data_out = 8'h85;
                    16'hABDB: data_out = 8'h86;
                    16'hABDC: data_out = 8'h87;
                    16'hABDD: data_out = 8'h88;
                    16'hABDE: data_out = 8'h89;
                    16'hABDF: data_out = 8'h8A;
                    16'hABE0: data_out = 8'h8B;
                    16'hABE1: data_out = 8'h8C;
                    16'hABE2: data_out = 8'h8D;
                    16'hABE3: data_out = 8'h8E;
                    16'hABE4: data_out = 8'h8F;
                    16'hABE5: data_out = 8'h90;
                    16'hABE6: data_out = 8'h91;
                    16'hABE7: data_out = 8'h92;
                    16'hABE8: data_out = 8'h93;
                    16'hABE9: data_out = 8'h94;
                    16'hABEA: data_out = 8'h95;
                    16'hABEB: data_out = 8'h96;
                    16'hABEC: data_out = 8'h97;
                    16'hABED: data_out = 8'h98;
                    16'hABEE: data_out = 8'h99;
                    16'hABEF: data_out = 8'h9A;
                    16'hABF0: data_out = 8'h9B;
                    16'hABF1: data_out = 8'h9C;
                    16'hABF2: data_out = 8'h9D;
                    16'hABF3: data_out = 8'h9E;
                    16'hABF4: data_out = 8'h9F;
                    16'hABF5: data_out = 8'hA0;
                    16'hABF6: data_out = 8'hA1;
                    16'hABF7: data_out = 8'hA2;
                    16'hABF8: data_out = 8'hA3;
                    16'hABF9: data_out = 8'hA4;
                    16'hABFA: data_out = 8'hA5;
                    16'hABFB: data_out = 8'hA6;
                    16'hABFC: data_out = 8'hA7;
                    16'hABFD: data_out = 8'hA8;
                    16'hABFE: data_out = 8'hA9;
                    16'hABFF: data_out = 8'hAA;
                    16'hAC00: data_out = 8'hAC;
                    16'hAC01: data_out = 8'hAB;
                    16'hAC02: data_out = 8'hAA;
                    16'hAC03: data_out = 8'hA9;
                    16'hAC04: data_out = 8'hA8;
                    16'hAC05: data_out = 8'hA7;
                    16'hAC06: data_out = 8'hA6;
                    16'hAC07: data_out = 8'hA5;
                    16'hAC08: data_out = 8'hA4;
                    16'hAC09: data_out = 8'hA3;
                    16'hAC0A: data_out = 8'hA2;
                    16'hAC0B: data_out = 8'hA1;
                    16'hAC0C: data_out = 8'hA0;
                    16'hAC0D: data_out = 8'h9F;
                    16'hAC0E: data_out = 8'h9E;
                    16'hAC0F: data_out = 8'h9D;
                    16'hAC10: data_out = 8'h9C;
                    16'hAC11: data_out = 8'h9B;
                    16'hAC12: data_out = 8'h9A;
                    16'hAC13: data_out = 8'h99;
                    16'hAC14: data_out = 8'h98;
                    16'hAC15: data_out = 8'h97;
                    16'hAC16: data_out = 8'h96;
                    16'hAC17: data_out = 8'h95;
                    16'hAC18: data_out = 8'h94;
                    16'hAC19: data_out = 8'h93;
                    16'hAC1A: data_out = 8'h92;
                    16'hAC1B: data_out = 8'h91;
                    16'hAC1C: data_out = 8'h90;
                    16'hAC1D: data_out = 8'h8F;
                    16'hAC1E: data_out = 8'h8E;
                    16'hAC1F: data_out = 8'h8D;
                    16'hAC20: data_out = 8'h8C;
                    16'hAC21: data_out = 8'h8B;
                    16'hAC22: data_out = 8'h8A;
                    16'hAC23: data_out = 8'h89;
                    16'hAC24: data_out = 8'h88;
                    16'hAC25: data_out = 8'h87;
                    16'hAC26: data_out = 8'h86;
                    16'hAC27: data_out = 8'h85;
                    16'hAC28: data_out = 8'h84;
                    16'hAC29: data_out = 8'h83;
                    16'hAC2A: data_out = 8'h82;
                    16'hAC2B: data_out = 8'h81;
                    16'hAC2C: data_out = 8'h0;
                    16'hAC2D: data_out = 8'h1;
                    16'hAC2E: data_out = 8'h2;
                    16'hAC2F: data_out = 8'h3;
                    16'hAC30: data_out = 8'h4;
                    16'hAC31: data_out = 8'h5;
                    16'hAC32: data_out = 8'h6;
                    16'hAC33: data_out = 8'h7;
                    16'hAC34: data_out = 8'h8;
                    16'hAC35: data_out = 8'h9;
                    16'hAC36: data_out = 8'hA;
                    16'hAC37: data_out = 8'hB;
                    16'hAC38: data_out = 8'hC;
                    16'hAC39: data_out = 8'hD;
                    16'hAC3A: data_out = 8'hE;
                    16'hAC3B: data_out = 8'hF;
                    16'hAC3C: data_out = 8'h10;
                    16'hAC3D: data_out = 8'h11;
                    16'hAC3E: data_out = 8'h12;
                    16'hAC3F: data_out = 8'h13;
                    16'hAC40: data_out = 8'h14;
                    16'hAC41: data_out = 8'h15;
                    16'hAC42: data_out = 8'h16;
                    16'hAC43: data_out = 8'h17;
                    16'hAC44: data_out = 8'h18;
                    16'hAC45: data_out = 8'h19;
                    16'hAC46: data_out = 8'h1A;
                    16'hAC47: data_out = 8'h1B;
                    16'hAC48: data_out = 8'h1C;
                    16'hAC49: data_out = 8'h1D;
                    16'hAC4A: data_out = 8'h1E;
                    16'hAC4B: data_out = 8'h1F;
                    16'hAC4C: data_out = 8'h20;
                    16'hAC4D: data_out = 8'h21;
                    16'hAC4E: data_out = 8'h22;
                    16'hAC4F: data_out = 8'h23;
                    16'hAC50: data_out = 8'h24;
                    16'hAC51: data_out = 8'h25;
                    16'hAC52: data_out = 8'h26;
                    16'hAC53: data_out = 8'h27;
                    16'hAC54: data_out = 8'h28;
                    16'hAC55: data_out = 8'h29;
                    16'hAC56: data_out = 8'h2A;
                    16'hAC57: data_out = 8'h2B;
                    16'hAC58: data_out = 8'h2C;
                    16'hAC59: data_out = 8'h2D;
                    16'hAC5A: data_out = 8'h2E;
                    16'hAC5B: data_out = 8'h2F;
                    16'hAC5C: data_out = 8'h30;
                    16'hAC5D: data_out = 8'h31;
                    16'hAC5E: data_out = 8'h32;
                    16'hAC5F: data_out = 8'h33;
                    16'hAC60: data_out = 8'h34;
                    16'hAC61: data_out = 8'h35;
                    16'hAC62: data_out = 8'h36;
                    16'hAC63: data_out = 8'h37;
                    16'hAC64: data_out = 8'h38;
                    16'hAC65: data_out = 8'h39;
                    16'hAC66: data_out = 8'h3A;
                    16'hAC67: data_out = 8'h3B;
                    16'hAC68: data_out = 8'h3C;
                    16'hAC69: data_out = 8'h3D;
                    16'hAC6A: data_out = 8'h3E;
                    16'hAC6B: data_out = 8'h3F;
                    16'hAC6C: data_out = 8'h40;
                    16'hAC6D: data_out = 8'h41;
                    16'hAC6E: data_out = 8'h42;
                    16'hAC6F: data_out = 8'h43;
                    16'hAC70: data_out = 8'h44;
                    16'hAC71: data_out = 8'h45;
                    16'hAC72: data_out = 8'h46;
                    16'hAC73: data_out = 8'h47;
                    16'hAC74: data_out = 8'h48;
                    16'hAC75: data_out = 8'h49;
                    16'hAC76: data_out = 8'h4A;
                    16'hAC77: data_out = 8'h4B;
                    16'hAC78: data_out = 8'h4C;
                    16'hAC79: data_out = 8'h4D;
                    16'hAC7A: data_out = 8'h4E;
                    16'hAC7B: data_out = 8'h4F;
                    16'hAC7C: data_out = 8'h50;
                    16'hAC7D: data_out = 8'h51;
                    16'hAC7E: data_out = 8'h52;
                    16'hAC7F: data_out = 8'h53;
                    16'hAC80: data_out = 8'hAC;
                    16'hAC81: data_out = 8'hAD;
                    16'hAC82: data_out = 8'hAE;
                    16'hAC83: data_out = 8'hAF;
                    16'hAC84: data_out = 8'hB0;
                    16'hAC85: data_out = 8'hB1;
                    16'hAC86: data_out = 8'hB2;
                    16'hAC87: data_out = 8'hB3;
                    16'hAC88: data_out = 8'hB4;
                    16'hAC89: data_out = 8'hB5;
                    16'hAC8A: data_out = 8'hB6;
                    16'hAC8B: data_out = 8'hB7;
                    16'hAC8C: data_out = 8'hB8;
                    16'hAC8D: data_out = 8'hB9;
                    16'hAC8E: data_out = 8'hBA;
                    16'hAC8F: data_out = 8'hBB;
                    16'hAC90: data_out = 8'hBC;
                    16'hAC91: data_out = 8'hBD;
                    16'hAC92: data_out = 8'hBE;
                    16'hAC93: data_out = 8'hBF;
                    16'hAC94: data_out = 8'hC0;
                    16'hAC95: data_out = 8'hC1;
                    16'hAC96: data_out = 8'hC2;
                    16'hAC97: data_out = 8'hC3;
                    16'hAC98: data_out = 8'hC4;
                    16'hAC99: data_out = 8'hC5;
                    16'hAC9A: data_out = 8'hC6;
                    16'hAC9B: data_out = 8'hC7;
                    16'hAC9C: data_out = 8'hC8;
                    16'hAC9D: data_out = 8'hC9;
                    16'hAC9E: data_out = 8'hCA;
                    16'hAC9F: data_out = 8'hCB;
                    16'hACA0: data_out = 8'hCC;
                    16'hACA1: data_out = 8'hCD;
                    16'hACA2: data_out = 8'hCE;
                    16'hACA3: data_out = 8'hCF;
                    16'hACA4: data_out = 8'hD0;
                    16'hACA5: data_out = 8'hD1;
                    16'hACA6: data_out = 8'hD2;
                    16'hACA7: data_out = 8'hD3;
                    16'hACA8: data_out = 8'hD4;
                    16'hACA9: data_out = 8'hD5;
                    16'hACAA: data_out = 8'hD6;
                    16'hACAB: data_out = 8'hD7;
                    16'hACAC: data_out = 8'hD8;
                    16'hACAD: data_out = 8'hD9;
                    16'hACAE: data_out = 8'hDA;
                    16'hACAF: data_out = 8'hDB;
                    16'hACB0: data_out = 8'hDC;
                    16'hACB1: data_out = 8'hDD;
                    16'hACB2: data_out = 8'hDE;
                    16'hACB3: data_out = 8'hDF;
                    16'hACB4: data_out = 8'hE0;
                    16'hACB5: data_out = 8'hE1;
                    16'hACB6: data_out = 8'hE2;
                    16'hACB7: data_out = 8'hE3;
                    16'hACB8: data_out = 8'hE4;
                    16'hACB9: data_out = 8'hE5;
                    16'hACBA: data_out = 8'hE6;
                    16'hACBB: data_out = 8'hE7;
                    16'hACBC: data_out = 8'hE8;
                    16'hACBD: data_out = 8'hE9;
                    16'hACBE: data_out = 8'hEA;
                    16'hACBF: data_out = 8'hEB;
                    16'hACC0: data_out = 8'hEC;
                    16'hACC1: data_out = 8'hED;
                    16'hACC2: data_out = 8'hEE;
                    16'hACC3: data_out = 8'hEF;
                    16'hACC4: data_out = 8'hF0;
                    16'hACC5: data_out = 8'hF1;
                    16'hACC6: data_out = 8'hF2;
                    16'hACC7: data_out = 8'hF3;
                    16'hACC8: data_out = 8'hF4;
                    16'hACC9: data_out = 8'hF5;
                    16'hACCA: data_out = 8'hF6;
                    16'hACCB: data_out = 8'hF7;
                    16'hACCC: data_out = 8'hF8;
                    16'hACCD: data_out = 8'hF9;
                    16'hACCE: data_out = 8'hFA;
                    16'hACCF: data_out = 8'hFB;
                    16'hACD0: data_out = 8'hFC;
                    16'hACD1: data_out = 8'hFD;
                    16'hACD2: data_out = 8'hFE;
                    16'hACD3: data_out = 8'hFF;
                    16'hACD4: data_out = 8'h80;
                    16'hACD5: data_out = 8'h81;
                    16'hACD6: data_out = 8'h82;
                    16'hACD7: data_out = 8'h83;
                    16'hACD8: data_out = 8'h84;
                    16'hACD9: data_out = 8'h85;
                    16'hACDA: data_out = 8'h86;
                    16'hACDB: data_out = 8'h87;
                    16'hACDC: data_out = 8'h88;
                    16'hACDD: data_out = 8'h89;
                    16'hACDE: data_out = 8'h8A;
                    16'hACDF: data_out = 8'h8B;
                    16'hACE0: data_out = 8'h8C;
                    16'hACE1: data_out = 8'h8D;
                    16'hACE2: data_out = 8'h8E;
                    16'hACE3: data_out = 8'h8F;
                    16'hACE4: data_out = 8'h90;
                    16'hACE5: data_out = 8'h91;
                    16'hACE6: data_out = 8'h92;
                    16'hACE7: data_out = 8'h93;
                    16'hACE8: data_out = 8'h94;
                    16'hACE9: data_out = 8'h95;
                    16'hACEA: data_out = 8'h96;
                    16'hACEB: data_out = 8'h97;
                    16'hACEC: data_out = 8'h98;
                    16'hACED: data_out = 8'h99;
                    16'hACEE: data_out = 8'h9A;
                    16'hACEF: data_out = 8'h9B;
                    16'hACF0: data_out = 8'h9C;
                    16'hACF1: data_out = 8'h9D;
                    16'hACF2: data_out = 8'h9E;
                    16'hACF3: data_out = 8'h9F;
                    16'hACF4: data_out = 8'hA0;
                    16'hACF5: data_out = 8'hA1;
                    16'hACF6: data_out = 8'hA2;
                    16'hACF7: data_out = 8'hA3;
                    16'hACF8: data_out = 8'hA4;
                    16'hACF9: data_out = 8'hA5;
                    16'hACFA: data_out = 8'hA6;
                    16'hACFB: data_out = 8'hA7;
                    16'hACFC: data_out = 8'hA8;
                    16'hACFD: data_out = 8'hA9;
                    16'hACFE: data_out = 8'hAA;
                    16'hACFF: data_out = 8'hAB;
                    16'hAD00: data_out = 8'hAD;
                    16'hAD01: data_out = 8'hAC;
                    16'hAD02: data_out = 8'hAB;
                    16'hAD03: data_out = 8'hAA;
                    16'hAD04: data_out = 8'hA9;
                    16'hAD05: data_out = 8'hA8;
                    16'hAD06: data_out = 8'hA7;
                    16'hAD07: data_out = 8'hA6;
                    16'hAD08: data_out = 8'hA5;
                    16'hAD09: data_out = 8'hA4;
                    16'hAD0A: data_out = 8'hA3;
                    16'hAD0B: data_out = 8'hA2;
                    16'hAD0C: data_out = 8'hA1;
                    16'hAD0D: data_out = 8'hA0;
                    16'hAD0E: data_out = 8'h9F;
                    16'hAD0F: data_out = 8'h9E;
                    16'hAD10: data_out = 8'h9D;
                    16'hAD11: data_out = 8'h9C;
                    16'hAD12: data_out = 8'h9B;
                    16'hAD13: data_out = 8'h9A;
                    16'hAD14: data_out = 8'h99;
                    16'hAD15: data_out = 8'h98;
                    16'hAD16: data_out = 8'h97;
                    16'hAD17: data_out = 8'h96;
                    16'hAD18: data_out = 8'h95;
                    16'hAD19: data_out = 8'h94;
                    16'hAD1A: data_out = 8'h93;
                    16'hAD1B: data_out = 8'h92;
                    16'hAD1C: data_out = 8'h91;
                    16'hAD1D: data_out = 8'h90;
                    16'hAD1E: data_out = 8'h8F;
                    16'hAD1F: data_out = 8'h8E;
                    16'hAD20: data_out = 8'h8D;
                    16'hAD21: data_out = 8'h8C;
                    16'hAD22: data_out = 8'h8B;
                    16'hAD23: data_out = 8'h8A;
                    16'hAD24: data_out = 8'h89;
                    16'hAD25: data_out = 8'h88;
                    16'hAD26: data_out = 8'h87;
                    16'hAD27: data_out = 8'h86;
                    16'hAD28: data_out = 8'h85;
                    16'hAD29: data_out = 8'h84;
                    16'hAD2A: data_out = 8'h83;
                    16'hAD2B: data_out = 8'h82;
                    16'hAD2C: data_out = 8'h81;
                    16'hAD2D: data_out = 8'h0;
                    16'hAD2E: data_out = 8'h1;
                    16'hAD2F: data_out = 8'h2;
                    16'hAD30: data_out = 8'h3;
                    16'hAD31: data_out = 8'h4;
                    16'hAD32: data_out = 8'h5;
                    16'hAD33: data_out = 8'h6;
                    16'hAD34: data_out = 8'h7;
                    16'hAD35: data_out = 8'h8;
                    16'hAD36: data_out = 8'h9;
                    16'hAD37: data_out = 8'hA;
                    16'hAD38: data_out = 8'hB;
                    16'hAD39: data_out = 8'hC;
                    16'hAD3A: data_out = 8'hD;
                    16'hAD3B: data_out = 8'hE;
                    16'hAD3C: data_out = 8'hF;
                    16'hAD3D: data_out = 8'h10;
                    16'hAD3E: data_out = 8'h11;
                    16'hAD3F: data_out = 8'h12;
                    16'hAD40: data_out = 8'h13;
                    16'hAD41: data_out = 8'h14;
                    16'hAD42: data_out = 8'h15;
                    16'hAD43: data_out = 8'h16;
                    16'hAD44: data_out = 8'h17;
                    16'hAD45: data_out = 8'h18;
                    16'hAD46: data_out = 8'h19;
                    16'hAD47: data_out = 8'h1A;
                    16'hAD48: data_out = 8'h1B;
                    16'hAD49: data_out = 8'h1C;
                    16'hAD4A: data_out = 8'h1D;
                    16'hAD4B: data_out = 8'h1E;
                    16'hAD4C: data_out = 8'h1F;
                    16'hAD4D: data_out = 8'h20;
                    16'hAD4E: data_out = 8'h21;
                    16'hAD4F: data_out = 8'h22;
                    16'hAD50: data_out = 8'h23;
                    16'hAD51: data_out = 8'h24;
                    16'hAD52: data_out = 8'h25;
                    16'hAD53: data_out = 8'h26;
                    16'hAD54: data_out = 8'h27;
                    16'hAD55: data_out = 8'h28;
                    16'hAD56: data_out = 8'h29;
                    16'hAD57: data_out = 8'h2A;
                    16'hAD58: data_out = 8'h2B;
                    16'hAD59: data_out = 8'h2C;
                    16'hAD5A: data_out = 8'h2D;
                    16'hAD5B: data_out = 8'h2E;
                    16'hAD5C: data_out = 8'h2F;
                    16'hAD5D: data_out = 8'h30;
                    16'hAD5E: data_out = 8'h31;
                    16'hAD5F: data_out = 8'h32;
                    16'hAD60: data_out = 8'h33;
                    16'hAD61: data_out = 8'h34;
                    16'hAD62: data_out = 8'h35;
                    16'hAD63: data_out = 8'h36;
                    16'hAD64: data_out = 8'h37;
                    16'hAD65: data_out = 8'h38;
                    16'hAD66: data_out = 8'h39;
                    16'hAD67: data_out = 8'h3A;
                    16'hAD68: data_out = 8'h3B;
                    16'hAD69: data_out = 8'h3C;
                    16'hAD6A: data_out = 8'h3D;
                    16'hAD6B: data_out = 8'h3E;
                    16'hAD6C: data_out = 8'h3F;
                    16'hAD6D: data_out = 8'h40;
                    16'hAD6E: data_out = 8'h41;
                    16'hAD6F: data_out = 8'h42;
                    16'hAD70: data_out = 8'h43;
                    16'hAD71: data_out = 8'h44;
                    16'hAD72: data_out = 8'h45;
                    16'hAD73: data_out = 8'h46;
                    16'hAD74: data_out = 8'h47;
                    16'hAD75: data_out = 8'h48;
                    16'hAD76: data_out = 8'h49;
                    16'hAD77: data_out = 8'h4A;
                    16'hAD78: data_out = 8'h4B;
                    16'hAD79: data_out = 8'h4C;
                    16'hAD7A: data_out = 8'h4D;
                    16'hAD7B: data_out = 8'h4E;
                    16'hAD7C: data_out = 8'h4F;
                    16'hAD7D: data_out = 8'h50;
                    16'hAD7E: data_out = 8'h51;
                    16'hAD7F: data_out = 8'h52;
                    16'hAD80: data_out = 8'hAD;
                    16'hAD81: data_out = 8'hAE;
                    16'hAD82: data_out = 8'hAF;
                    16'hAD83: data_out = 8'hB0;
                    16'hAD84: data_out = 8'hB1;
                    16'hAD85: data_out = 8'hB2;
                    16'hAD86: data_out = 8'hB3;
                    16'hAD87: data_out = 8'hB4;
                    16'hAD88: data_out = 8'hB5;
                    16'hAD89: data_out = 8'hB6;
                    16'hAD8A: data_out = 8'hB7;
                    16'hAD8B: data_out = 8'hB8;
                    16'hAD8C: data_out = 8'hB9;
                    16'hAD8D: data_out = 8'hBA;
                    16'hAD8E: data_out = 8'hBB;
                    16'hAD8F: data_out = 8'hBC;
                    16'hAD90: data_out = 8'hBD;
                    16'hAD91: data_out = 8'hBE;
                    16'hAD92: data_out = 8'hBF;
                    16'hAD93: data_out = 8'hC0;
                    16'hAD94: data_out = 8'hC1;
                    16'hAD95: data_out = 8'hC2;
                    16'hAD96: data_out = 8'hC3;
                    16'hAD97: data_out = 8'hC4;
                    16'hAD98: data_out = 8'hC5;
                    16'hAD99: data_out = 8'hC6;
                    16'hAD9A: data_out = 8'hC7;
                    16'hAD9B: data_out = 8'hC8;
                    16'hAD9C: data_out = 8'hC9;
                    16'hAD9D: data_out = 8'hCA;
                    16'hAD9E: data_out = 8'hCB;
                    16'hAD9F: data_out = 8'hCC;
                    16'hADA0: data_out = 8'hCD;
                    16'hADA1: data_out = 8'hCE;
                    16'hADA2: data_out = 8'hCF;
                    16'hADA3: data_out = 8'hD0;
                    16'hADA4: data_out = 8'hD1;
                    16'hADA5: data_out = 8'hD2;
                    16'hADA6: data_out = 8'hD3;
                    16'hADA7: data_out = 8'hD4;
                    16'hADA8: data_out = 8'hD5;
                    16'hADA9: data_out = 8'hD6;
                    16'hADAA: data_out = 8'hD7;
                    16'hADAB: data_out = 8'hD8;
                    16'hADAC: data_out = 8'hD9;
                    16'hADAD: data_out = 8'hDA;
                    16'hADAE: data_out = 8'hDB;
                    16'hADAF: data_out = 8'hDC;
                    16'hADB0: data_out = 8'hDD;
                    16'hADB1: data_out = 8'hDE;
                    16'hADB2: data_out = 8'hDF;
                    16'hADB3: data_out = 8'hE0;
                    16'hADB4: data_out = 8'hE1;
                    16'hADB5: data_out = 8'hE2;
                    16'hADB6: data_out = 8'hE3;
                    16'hADB7: data_out = 8'hE4;
                    16'hADB8: data_out = 8'hE5;
                    16'hADB9: data_out = 8'hE6;
                    16'hADBA: data_out = 8'hE7;
                    16'hADBB: data_out = 8'hE8;
                    16'hADBC: data_out = 8'hE9;
                    16'hADBD: data_out = 8'hEA;
                    16'hADBE: data_out = 8'hEB;
                    16'hADBF: data_out = 8'hEC;
                    16'hADC0: data_out = 8'hED;
                    16'hADC1: data_out = 8'hEE;
                    16'hADC2: data_out = 8'hEF;
                    16'hADC3: data_out = 8'hF0;
                    16'hADC4: data_out = 8'hF1;
                    16'hADC5: data_out = 8'hF2;
                    16'hADC6: data_out = 8'hF3;
                    16'hADC7: data_out = 8'hF4;
                    16'hADC8: data_out = 8'hF5;
                    16'hADC9: data_out = 8'hF6;
                    16'hADCA: data_out = 8'hF7;
                    16'hADCB: data_out = 8'hF8;
                    16'hADCC: data_out = 8'hF9;
                    16'hADCD: data_out = 8'hFA;
                    16'hADCE: data_out = 8'hFB;
                    16'hADCF: data_out = 8'hFC;
                    16'hADD0: data_out = 8'hFD;
                    16'hADD1: data_out = 8'hFE;
                    16'hADD2: data_out = 8'hFF;
                    16'hADD3: data_out = 8'h80;
                    16'hADD4: data_out = 8'h81;
                    16'hADD5: data_out = 8'h82;
                    16'hADD6: data_out = 8'h83;
                    16'hADD7: data_out = 8'h84;
                    16'hADD8: data_out = 8'h85;
                    16'hADD9: data_out = 8'h86;
                    16'hADDA: data_out = 8'h87;
                    16'hADDB: data_out = 8'h88;
                    16'hADDC: data_out = 8'h89;
                    16'hADDD: data_out = 8'h8A;
                    16'hADDE: data_out = 8'h8B;
                    16'hADDF: data_out = 8'h8C;
                    16'hADE0: data_out = 8'h8D;
                    16'hADE1: data_out = 8'h8E;
                    16'hADE2: data_out = 8'h8F;
                    16'hADE3: data_out = 8'h90;
                    16'hADE4: data_out = 8'h91;
                    16'hADE5: data_out = 8'h92;
                    16'hADE6: data_out = 8'h93;
                    16'hADE7: data_out = 8'h94;
                    16'hADE8: data_out = 8'h95;
                    16'hADE9: data_out = 8'h96;
                    16'hADEA: data_out = 8'h97;
                    16'hADEB: data_out = 8'h98;
                    16'hADEC: data_out = 8'h99;
                    16'hADED: data_out = 8'h9A;
                    16'hADEE: data_out = 8'h9B;
                    16'hADEF: data_out = 8'h9C;
                    16'hADF0: data_out = 8'h9D;
                    16'hADF1: data_out = 8'h9E;
                    16'hADF2: data_out = 8'h9F;
                    16'hADF3: data_out = 8'hA0;
                    16'hADF4: data_out = 8'hA1;
                    16'hADF5: data_out = 8'hA2;
                    16'hADF6: data_out = 8'hA3;
                    16'hADF7: data_out = 8'hA4;
                    16'hADF8: data_out = 8'hA5;
                    16'hADF9: data_out = 8'hA6;
                    16'hADFA: data_out = 8'hA7;
                    16'hADFB: data_out = 8'hA8;
                    16'hADFC: data_out = 8'hA9;
                    16'hADFD: data_out = 8'hAA;
                    16'hADFE: data_out = 8'hAB;
                    16'hADFF: data_out = 8'hAC;
                    16'hAE00: data_out = 8'hAE;
                    16'hAE01: data_out = 8'hAD;
                    16'hAE02: data_out = 8'hAC;
                    16'hAE03: data_out = 8'hAB;
                    16'hAE04: data_out = 8'hAA;
                    16'hAE05: data_out = 8'hA9;
                    16'hAE06: data_out = 8'hA8;
                    16'hAE07: data_out = 8'hA7;
                    16'hAE08: data_out = 8'hA6;
                    16'hAE09: data_out = 8'hA5;
                    16'hAE0A: data_out = 8'hA4;
                    16'hAE0B: data_out = 8'hA3;
                    16'hAE0C: data_out = 8'hA2;
                    16'hAE0D: data_out = 8'hA1;
                    16'hAE0E: data_out = 8'hA0;
                    16'hAE0F: data_out = 8'h9F;
                    16'hAE10: data_out = 8'h9E;
                    16'hAE11: data_out = 8'h9D;
                    16'hAE12: data_out = 8'h9C;
                    16'hAE13: data_out = 8'h9B;
                    16'hAE14: data_out = 8'h9A;
                    16'hAE15: data_out = 8'h99;
                    16'hAE16: data_out = 8'h98;
                    16'hAE17: data_out = 8'h97;
                    16'hAE18: data_out = 8'h96;
                    16'hAE19: data_out = 8'h95;
                    16'hAE1A: data_out = 8'h94;
                    16'hAE1B: data_out = 8'h93;
                    16'hAE1C: data_out = 8'h92;
                    16'hAE1D: data_out = 8'h91;
                    16'hAE1E: data_out = 8'h90;
                    16'hAE1F: data_out = 8'h8F;
                    16'hAE20: data_out = 8'h8E;
                    16'hAE21: data_out = 8'h8D;
                    16'hAE22: data_out = 8'h8C;
                    16'hAE23: data_out = 8'h8B;
                    16'hAE24: data_out = 8'h8A;
                    16'hAE25: data_out = 8'h89;
                    16'hAE26: data_out = 8'h88;
                    16'hAE27: data_out = 8'h87;
                    16'hAE28: data_out = 8'h86;
                    16'hAE29: data_out = 8'h85;
                    16'hAE2A: data_out = 8'h84;
                    16'hAE2B: data_out = 8'h83;
                    16'hAE2C: data_out = 8'h82;
                    16'hAE2D: data_out = 8'h81;
                    16'hAE2E: data_out = 8'h0;
                    16'hAE2F: data_out = 8'h1;
                    16'hAE30: data_out = 8'h2;
                    16'hAE31: data_out = 8'h3;
                    16'hAE32: data_out = 8'h4;
                    16'hAE33: data_out = 8'h5;
                    16'hAE34: data_out = 8'h6;
                    16'hAE35: data_out = 8'h7;
                    16'hAE36: data_out = 8'h8;
                    16'hAE37: data_out = 8'h9;
                    16'hAE38: data_out = 8'hA;
                    16'hAE39: data_out = 8'hB;
                    16'hAE3A: data_out = 8'hC;
                    16'hAE3B: data_out = 8'hD;
                    16'hAE3C: data_out = 8'hE;
                    16'hAE3D: data_out = 8'hF;
                    16'hAE3E: data_out = 8'h10;
                    16'hAE3F: data_out = 8'h11;
                    16'hAE40: data_out = 8'h12;
                    16'hAE41: data_out = 8'h13;
                    16'hAE42: data_out = 8'h14;
                    16'hAE43: data_out = 8'h15;
                    16'hAE44: data_out = 8'h16;
                    16'hAE45: data_out = 8'h17;
                    16'hAE46: data_out = 8'h18;
                    16'hAE47: data_out = 8'h19;
                    16'hAE48: data_out = 8'h1A;
                    16'hAE49: data_out = 8'h1B;
                    16'hAE4A: data_out = 8'h1C;
                    16'hAE4B: data_out = 8'h1D;
                    16'hAE4C: data_out = 8'h1E;
                    16'hAE4D: data_out = 8'h1F;
                    16'hAE4E: data_out = 8'h20;
                    16'hAE4F: data_out = 8'h21;
                    16'hAE50: data_out = 8'h22;
                    16'hAE51: data_out = 8'h23;
                    16'hAE52: data_out = 8'h24;
                    16'hAE53: data_out = 8'h25;
                    16'hAE54: data_out = 8'h26;
                    16'hAE55: data_out = 8'h27;
                    16'hAE56: data_out = 8'h28;
                    16'hAE57: data_out = 8'h29;
                    16'hAE58: data_out = 8'h2A;
                    16'hAE59: data_out = 8'h2B;
                    16'hAE5A: data_out = 8'h2C;
                    16'hAE5B: data_out = 8'h2D;
                    16'hAE5C: data_out = 8'h2E;
                    16'hAE5D: data_out = 8'h2F;
                    16'hAE5E: data_out = 8'h30;
                    16'hAE5F: data_out = 8'h31;
                    16'hAE60: data_out = 8'h32;
                    16'hAE61: data_out = 8'h33;
                    16'hAE62: data_out = 8'h34;
                    16'hAE63: data_out = 8'h35;
                    16'hAE64: data_out = 8'h36;
                    16'hAE65: data_out = 8'h37;
                    16'hAE66: data_out = 8'h38;
                    16'hAE67: data_out = 8'h39;
                    16'hAE68: data_out = 8'h3A;
                    16'hAE69: data_out = 8'h3B;
                    16'hAE6A: data_out = 8'h3C;
                    16'hAE6B: data_out = 8'h3D;
                    16'hAE6C: data_out = 8'h3E;
                    16'hAE6D: data_out = 8'h3F;
                    16'hAE6E: data_out = 8'h40;
                    16'hAE6F: data_out = 8'h41;
                    16'hAE70: data_out = 8'h42;
                    16'hAE71: data_out = 8'h43;
                    16'hAE72: data_out = 8'h44;
                    16'hAE73: data_out = 8'h45;
                    16'hAE74: data_out = 8'h46;
                    16'hAE75: data_out = 8'h47;
                    16'hAE76: data_out = 8'h48;
                    16'hAE77: data_out = 8'h49;
                    16'hAE78: data_out = 8'h4A;
                    16'hAE79: data_out = 8'h4B;
                    16'hAE7A: data_out = 8'h4C;
                    16'hAE7B: data_out = 8'h4D;
                    16'hAE7C: data_out = 8'h4E;
                    16'hAE7D: data_out = 8'h4F;
                    16'hAE7E: data_out = 8'h50;
                    16'hAE7F: data_out = 8'h51;
                    16'hAE80: data_out = 8'hAE;
                    16'hAE81: data_out = 8'hAF;
                    16'hAE82: data_out = 8'hB0;
                    16'hAE83: data_out = 8'hB1;
                    16'hAE84: data_out = 8'hB2;
                    16'hAE85: data_out = 8'hB3;
                    16'hAE86: data_out = 8'hB4;
                    16'hAE87: data_out = 8'hB5;
                    16'hAE88: data_out = 8'hB6;
                    16'hAE89: data_out = 8'hB7;
                    16'hAE8A: data_out = 8'hB8;
                    16'hAE8B: data_out = 8'hB9;
                    16'hAE8C: data_out = 8'hBA;
                    16'hAE8D: data_out = 8'hBB;
                    16'hAE8E: data_out = 8'hBC;
                    16'hAE8F: data_out = 8'hBD;
                    16'hAE90: data_out = 8'hBE;
                    16'hAE91: data_out = 8'hBF;
                    16'hAE92: data_out = 8'hC0;
                    16'hAE93: data_out = 8'hC1;
                    16'hAE94: data_out = 8'hC2;
                    16'hAE95: data_out = 8'hC3;
                    16'hAE96: data_out = 8'hC4;
                    16'hAE97: data_out = 8'hC5;
                    16'hAE98: data_out = 8'hC6;
                    16'hAE99: data_out = 8'hC7;
                    16'hAE9A: data_out = 8'hC8;
                    16'hAE9B: data_out = 8'hC9;
                    16'hAE9C: data_out = 8'hCA;
                    16'hAE9D: data_out = 8'hCB;
                    16'hAE9E: data_out = 8'hCC;
                    16'hAE9F: data_out = 8'hCD;
                    16'hAEA0: data_out = 8'hCE;
                    16'hAEA1: data_out = 8'hCF;
                    16'hAEA2: data_out = 8'hD0;
                    16'hAEA3: data_out = 8'hD1;
                    16'hAEA4: data_out = 8'hD2;
                    16'hAEA5: data_out = 8'hD3;
                    16'hAEA6: data_out = 8'hD4;
                    16'hAEA7: data_out = 8'hD5;
                    16'hAEA8: data_out = 8'hD6;
                    16'hAEA9: data_out = 8'hD7;
                    16'hAEAA: data_out = 8'hD8;
                    16'hAEAB: data_out = 8'hD9;
                    16'hAEAC: data_out = 8'hDA;
                    16'hAEAD: data_out = 8'hDB;
                    16'hAEAE: data_out = 8'hDC;
                    16'hAEAF: data_out = 8'hDD;
                    16'hAEB0: data_out = 8'hDE;
                    16'hAEB1: data_out = 8'hDF;
                    16'hAEB2: data_out = 8'hE0;
                    16'hAEB3: data_out = 8'hE1;
                    16'hAEB4: data_out = 8'hE2;
                    16'hAEB5: data_out = 8'hE3;
                    16'hAEB6: data_out = 8'hE4;
                    16'hAEB7: data_out = 8'hE5;
                    16'hAEB8: data_out = 8'hE6;
                    16'hAEB9: data_out = 8'hE7;
                    16'hAEBA: data_out = 8'hE8;
                    16'hAEBB: data_out = 8'hE9;
                    16'hAEBC: data_out = 8'hEA;
                    16'hAEBD: data_out = 8'hEB;
                    16'hAEBE: data_out = 8'hEC;
                    16'hAEBF: data_out = 8'hED;
                    16'hAEC0: data_out = 8'hEE;
                    16'hAEC1: data_out = 8'hEF;
                    16'hAEC2: data_out = 8'hF0;
                    16'hAEC3: data_out = 8'hF1;
                    16'hAEC4: data_out = 8'hF2;
                    16'hAEC5: data_out = 8'hF3;
                    16'hAEC6: data_out = 8'hF4;
                    16'hAEC7: data_out = 8'hF5;
                    16'hAEC8: data_out = 8'hF6;
                    16'hAEC9: data_out = 8'hF7;
                    16'hAECA: data_out = 8'hF8;
                    16'hAECB: data_out = 8'hF9;
                    16'hAECC: data_out = 8'hFA;
                    16'hAECD: data_out = 8'hFB;
                    16'hAECE: data_out = 8'hFC;
                    16'hAECF: data_out = 8'hFD;
                    16'hAED0: data_out = 8'hFE;
                    16'hAED1: data_out = 8'hFF;
                    16'hAED2: data_out = 8'h80;
                    16'hAED3: data_out = 8'h81;
                    16'hAED4: data_out = 8'h82;
                    16'hAED5: data_out = 8'h83;
                    16'hAED6: data_out = 8'h84;
                    16'hAED7: data_out = 8'h85;
                    16'hAED8: data_out = 8'h86;
                    16'hAED9: data_out = 8'h87;
                    16'hAEDA: data_out = 8'h88;
                    16'hAEDB: data_out = 8'h89;
                    16'hAEDC: data_out = 8'h8A;
                    16'hAEDD: data_out = 8'h8B;
                    16'hAEDE: data_out = 8'h8C;
                    16'hAEDF: data_out = 8'h8D;
                    16'hAEE0: data_out = 8'h8E;
                    16'hAEE1: data_out = 8'h8F;
                    16'hAEE2: data_out = 8'h90;
                    16'hAEE3: data_out = 8'h91;
                    16'hAEE4: data_out = 8'h92;
                    16'hAEE5: data_out = 8'h93;
                    16'hAEE6: data_out = 8'h94;
                    16'hAEE7: data_out = 8'h95;
                    16'hAEE8: data_out = 8'h96;
                    16'hAEE9: data_out = 8'h97;
                    16'hAEEA: data_out = 8'h98;
                    16'hAEEB: data_out = 8'h99;
                    16'hAEEC: data_out = 8'h9A;
                    16'hAEED: data_out = 8'h9B;
                    16'hAEEE: data_out = 8'h9C;
                    16'hAEEF: data_out = 8'h9D;
                    16'hAEF0: data_out = 8'h9E;
                    16'hAEF1: data_out = 8'h9F;
                    16'hAEF2: data_out = 8'hA0;
                    16'hAEF3: data_out = 8'hA1;
                    16'hAEF4: data_out = 8'hA2;
                    16'hAEF5: data_out = 8'hA3;
                    16'hAEF6: data_out = 8'hA4;
                    16'hAEF7: data_out = 8'hA5;
                    16'hAEF8: data_out = 8'hA6;
                    16'hAEF9: data_out = 8'hA7;
                    16'hAEFA: data_out = 8'hA8;
                    16'hAEFB: data_out = 8'hA9;
                    16'hAEFC: data_out = 8'hAA;
                    16'hAEFD: data_out = 8'hAB;
                    16'hAEFE: data_out = 8'hAC;
                    16'hAEFF: data_out = 8'hAD;
                    16'hAF00: data_out = 8'hAF;
                    16'hAF01: data_out = 8'hAE;
                    16'hAF02: data_out = 8'hAD;
                    16'hAF03: data_out = 8'hAC;
                    16'hAF04: data_out = 8'hAB;
                    16'hAF05: data_out = 8'hAA;
                    16'hAF06: data_out = 8'hA9;
                    16'hAF07: data_out = 8'hA8;
                    16'hAF08: data_out = 8'hA7;
                    16'hAF09: data_out = 8'hA6;
                    16'hAF0A: data_out = 8'hA5;
                    16'hAF0B: data_out = 8'hA4;
                    16'hAF0C: data_out = 8'hA3;
                    16'hAF0D: data_out = 8'hA2;
                    16'hAF0E: data_out = 8'hA1;
                    16'hAF0F: data_out = 8'hA0;
                    16'hAF10: data_out = 8'h9F;
                    16'hAF11: data_out = 8'h9E;
                    16'hAF12: data_out = 8'h9D;
                    16'hAF13: data_out = 8'h9C;
                    16'hAF14: data_out = 8'h9B;
                    16'hAF15: data_out = 8'h9A;
                    16'hAF16: data_out = 8'h99;
                    16'hAF17: data_out = 8'h98;
                    16'hAF18: data_out = 8'h97;
                    16'hAF19: data_out = 8'h96;
                    16'hAF1A: data_out = 8'h95;
                    16'hAF1B: data_out = 8'h94;
                    16'hAF1C: data_out = 8'h93;
                    16'hAF1D: data_out = 8'h92;
                    16'hAF1E: data_out = 8'h91;
                    16'hAF1F: data_out = 8'h90;
                    16'hAF20: data_out = 8'h8F;
                    16'hAF21: data_out = 8'h8E;
                    16'hAF22: data_out = 8'h8D;
                    16'hAF23: data_out = 8'h8C;
                    16'hAF24: data_out = 8'h8B;
                    16'hAF25: data_out = 8'h8A;
                    16'hAF26: data_out = 8'h89;
                    16'hAF27: data_out = 8'h88;
                    16'hAF28: data_out = 8'h87;
                    16'hAF29: data_out = 8'h86;
                    16'hAF2A: data_out = 8'h85;
                    16'hAF2B: data_out = 8'h84;
                    16'hAF2C: data_out = 8'h83;
                    16'hAF2D: data_out = 8'h82;
                    16'hAF2E: data_out = 8'h81;
                    16'hAF2F: data_out = 8'h0;
                    16'hAF30: data_out = 8'h1;
                    16'hAF31: data_out = 8'h2;
                    16'hAF32: data_out = 8'h3;
                    16'hAF33: data_out = 8'h4;
                    16'hAF34: data_out = 8'h5;
                    16'hAF35: data_out = 8'h6;
                    16'hAF36: data_out = 8'h7;
                    16'hAF37: data_out = 8'h8;
                    16'hAF38: data_out = 8'h9;
                    16'hAF39: data_out = 8'hA;
                    16'hAF3A: data_out = 8'hB;
                    16'hAF3B: data_out = 8'hC;
                    16'hAF3C: data_out = 8'hD;
                    16'hAF3D: data_out = 8'hE;
                    16'hAF3E: data_out = 8'hF;
                    16'hAF3F: data_out = 8'h10;
                    16'hAF40: data_out = 8'h11;
                    16'hAF41: data_out = 8'h12;
                    16'hAF42: data_out = 8'h13;
                    16'hAF43: data_out = 8'h14;
                    16'hAF44: data_out = 8'h15;
                    16'hAF45: data_out = 8'h16;
                    16'hAF46: data_out = 8'h17;
                    16'hAF47: data_out = 8'h18;
                    16'hAF48: data_out = 8'h19;
                    16'hAF49: data_out = 8'h1A;
                    16'hAF4A: data_out = 8'h1B;
                    16'hAF4B: data_out = 8'h1C;
                    16'hAF4C: data_out = 8'h1D;
                    16'hAF4D: data_out = 8'h1E;
                    16'hAF4E: data_out = 8'h1F;
                    16'hAF4F: data_out = 8'h20;
                    16'hAF50: data_out = 8'h21;
                    16'hAF51: data_out = 8'h22;
                    16'hAF52: data_out = 8'h23;
                    16'hAF53: data_out = 8'h24;
                    16'hAF54: data_out = 8'h25;
                    16'hAF55: data_out = 8'h26;
                    16'hAF56: data_out = 8'h27;
                    16'hAF57: data_out = 8'h28;
                    16'hAF58: data_out = 8'h29;
                    16'hAF59: data_out = 8'h2A;
                    16'hAF5A: data_out = 8'h2B;
                    16'hAF5B: data_out = 8'h2C;
                    16'hAF5C: data_out = 8'h2D;
                    16'hAF5D: data_out = 8'h2E;
                    16'hAF5E: data_out = 8'h2F;
                    16'hAF5F: data_out = 8'h30;
                    16'hAF60: data_out = 8'h31;
                    16'hAF61: data_out = 8'h32;
                    16'hAF62: data_out = 8'h33;
                    16'hAF63: data_out = 8'h34;
                    16'hAF64: data_out = 8'h35;
                    16'hAF65: data_out = 8'h36;
                    16'hAF66: data_out = 8'h37;
                    16'hAF67: data_out = 8'h38;
                    16'hAF68: data_out = 8'h39;
                    16'hAF69: data_out = 8'h3A;
                    16'hAF6A: data_out = 8'h3B;
                    16'hAF6B: data_out = 8'h3C;
                    16'hAF6C: data_out = 8'h3D;
                    16'hAF6D: data_out = 8'h3E;
                    16'hAF6E: data_out = 8'h3F;
                    16'hAF6F: data_out = 8'h40;
                    16'hAF70: data_out = 8'h41;
                    16'hAF71: data_out = 8'h42;
                    16'hAF72: data_out = 8'h43;
                    16'hAF73: data_out = 8'h44;
                    16'hAF74: data_out = 8'h45;
                    16'hAF75: data_out = 8'h46;
                    16'hAF76: data_out = 8'h47;
                    16'hAF77: data_out = 8'h48;
                    16'hAF78: data_out = 8'h49;
                    16'hAF79: data_out = 8'h4A;
                    16'hAF7A: data_out = 8'h4B;
                    16'hAF7B: data_out = 8'h4C;
                    16'hAF7C: data_out = 8'h4D;
                    16'hAF7D: data_out = 8'h4E;
                    16'hAF7E: data_out = 8'h4F;
                    16'hAF7F: data_out = 8'h50;
                    16'hAF80: data_out = 8'hAF;
                    16'hAF81: data_out = 8'hB0;
                    16'hAF82: data_out = 8'hB1;
                    16'hAF83: data_out = 8'hB2;
                    16'hAF84: data_out = 8'hB3;
                    16'hAF85: data_out = 8'hB4;
                    16'hAF86: data_out = 8'hB5;
                    16'hAF87: data_out = 8'hB6;
                    16'hAF88: data_out = 8'hB7;
                    16'hAF89: data_out = 8'hB8;
                    16'hAF8A: data_out = 8'hB9;
                    16'hAF8B: data_out = 8'hBA;
                    16'hAF8C: data_out = 8'hBB;
                    16'hAF8D: data_out = 8'hBC;
                    16'hAF8E: data_out = 8'hBD;
                    16'hAF8F: data_out = 8'hBE;
                    16'hAF90: data_out = 8'hBF;
                    16'hAF91: data_out = 8'hC0;
                    16'hAF92: data_out = 8'hC1;
                    16'hAF93: data_out = 8'hC2;
                    16'hAF94: data_out = 8'hC3;
                    16'hAF95: data_out = 8'hC4;
                    16'hAF96: data_out = 8'hC5;
                    16'hAF97: data_out = 8'hC6;
                    16'hAF98: data_out = 8'hC7;
                    16'hAF99: data_out = 8'hC8;
                    16'hAF9A: data_out = 8'hC9;
                    16'hAF9B: data_out = 8'hCA;
                    16'hAF9C: data_out = 8'hCB;
                    16'hAF9D: data_out = 8'hCC;
                    16'hAF9E: data_out = 8'hCD;
                    16'hAF9F: data_out = 8'hCE;
                    16'hAFA0: data_out = 8'hCF;
                    16'hAFA1: data_out = 8'hD0;
                    16'hAFA2: data_out = 8'hD1;
                    16'hAFA3: data_out = 8'hD2;
                    16'hAFA4: data_out = 8'hD3;
                    16'hAFA5: data_out = 8'hD4;
                    16'hAFA6: data_out = 8'hD5;
                    16'hAFA7: data_out = 8'hD6;
                    16'hAFA8: data_out = 8'hD7;
                    16'hAFA9: data_out = 8'hD8;
                    16'hAFAA: data_out = 8'hD9;
                    16'hAFAB: data_out = 8'hDA;
                    16'hAFAC: data_out = 8'hDB;
                    16'hAFAD: data_out = 8'hDC;
                    16'hAFAE: data_out = 8'hDD;
                    16'hAFAF: data_out = 8'hDE;
                    16'hAFB0: data_out = 8'hDF;
                    16'hAFB1: data_out = 8'hE0;
                    16'hAFB2: data_out = 8'hE1;
                    16'hAFB3: data_out = 8'hE2;
                    16'hAFB4: data_out = 8'hE3;
                    16'hAFB5: data_out = 8'hE4;
                    16'hAFB6: data_out = 8'hE5;
                    16'hAFB7: data_out = 8'hE6;
                    16'hAFB8: data_out = 8'hE7;
                    16'hAFB9: data_out = 8'hE8;
                    16'hAFBA: data_out = 8'hE9;
                    16'hAFBB: data_out = 8'hEA;
                    16'hAFBC: data_out = 8'hEB;
                    16'hAFBD: data_out = 8'hEC;
                    16'hAFBE: data_out = 8'hED;
                    16'hAFBF: data_out = 8'hEE;
                    16'hAFC0: data_out = 8'hEF;
                    16'hAFC1: data_out = 8'hF0;
                    16'hAFC2: data_out = 8'hF1;
                    16'hAFC3: data_out = 8'hF2;
                    16'hAFC4: data_out = 8'hF3;
                    16'hAFC5: data_out = 8'hF4;
                    16'hAFC6: data_out = 8'hF5;
                    16'hAFC7: data_out = 8'hF6;
                    16'hAFC8: data_out = 8'hF7;
                    16'hAFC9: data_out = 8'hF8;
                    16'hAFCA: data_out = 8'hF9;
                    16'hAFCB: data_out = 8'hFA;
                    16'hAFCC: data_out = 8'hFB;
                    16'hAFCD: data_out = 8'hFC;
                    16'hAFCE: data_out = 8'hFD;
                    16'hAFCF: data_out = 8'hFE;
                    16'hAFD0: data_out = 8'hFF;
                    16'hAFD1: data_out = 8'h80;
                    16'hAFD2: data_out = 8'h81;
                    16'hAFD3: data_out = 8'h82;
                    16'hAFD4: data_out = 8'h83;
                    16'hAFD5: data_out = 8'h84;
                    16'hAFD6: data_out = 8'h85;
                    16'hAFD7: data_out = 8'h86;
                    16'hAFD8: data_out = 8'h87;
                    16'hAFD9: data_out = 8'h88;
                    16'hAFDA: data_out = 8'h89;
                    16'hAFDB: data_out = 8'h8A;
                    16'hAFDC: data_out = 8'h8B;
                    16'hAFDD: data_out = 8'h8C;
                    16'hAFDE: data_out = 8'h8D;
                    16'hAFDF: data_out = 8'h8E;
                    16'hAFE0: data_out = 8'h8F;
                    16'hAFE1: data_out = 8'h90;
                    16'hAFE2: data_out = 8'h91;
                    16'hAFE3: data_out = 8'h92;
                    16'hAFE4: data_out = 8'h93;
                    16'hAFE5: data_out = 8'h94;
                    16'hAFE6: data_out = 8'h95;
                    16'hAFE7: data_out = 8'h96;
                    16'hAFE8: data_out = 8'h97;
                    16'hAFE9: data_out = 8'h98;
                    16'hAFEA: data_out = 8'h99;
                    16'hAFEB: data_out = 8'h9A;
                    16'hAFEC: data_out = 8'h9B;
                    16'hAFED: data_out = 8'h9C;
                    16'hAFEE: data_out = 8'h9D;
                    16'hAFEF: data_out = 8'h9E;
                    16'hAFF0: data_out = 8'h9F;
                    16'hAFF1: data_out = 8'hA0;
                    16'hAFF2: data_out = 8'hA1;
                    16'hAFF3: data_out = 8'hA2;
                    16'hAFF4: data_out = 8'hA3;
                    16'hAFF5: data_out = 8'hA4;
                    16'hAFF6: data_out = 8'hA5;
                    16'hAFF7: data_out = 8'hA6;
                    16'hAFF8: data_out = 8'hA7;
                    16'hAFF9: data_out = 8'hA8;
                    16'hAFFA: data_out = 8'hA9;
                    16'hAFFB: data_out = 8'hAA;
                    16'hAFFC: data_out = 8'hAB;
                    16'hAFFD: data_out = 8'hAC;
                    16'hAFFE: data_out = 8'hAD;
                    16'hAFFF: data_out = 8'hAE;
                    16'hB000: data_out = 8'hB0;
                    16'hB001: data_out = 8'hAF;
                    16'hB002: data_out = 8'hAE;
                    16'hB003: data_out = 8'hAD;
                    16'hB004: data_out = 8'hAC;
                    16'hB005: data_out = 8'hAB;
                    16'hB006: data_out = 8'hAA;
                    16'hB007: data_out = 8'hA9;
                    16'hB008: data_out = 8'hA8;
                    16'hB009: data_out = 8'hA7;
                    16'hB00A: data_out = 8'hA6;
                    16'hB00B: data_out = 8'hA5;
                    16'hB00C: data_out = 8'hA4;
                    16'hB00D: data_out = 8'hA3;
                    16'hB00E: data_out = 8'hA2;
                    16'hB00F: data_out = 8'hA1;
                    16'hB010: data_out = 8'hA0;
                    16'hB011: data_out = 8'h9F;
                    16'hB012: data_out = 8'h9E;
                    16'hB013: data_out = 8'h9D;
                    16'hB014: data_out = 8'h9C;
                    16'hB015: data_out = 8'h9B;
                    16'hB016: data_out = 8'h9A;
                    16'hB017: data_out = 8'h99;
                    16'hB018: data_out = 8'h98;
                    16'hB019: data_out = 8'h97;
                    16'hB01A: data_out = 8'h96;
                    16'hB01B: data_out = 8'h95;
                    16'hB01C: data_out = 8'h94;
                    16'hB01D: data_out = 8'h93;
                    16'hB01E: data_out = 8'h92;
                    16'hB01F: data_out = 8'h91;
                    16'hB020: data_out = 8'h90;
                    16'hB021: data_out = 8'h8F;
                    16'hB022: data_out = 8'h8E;
                    16'hB023: data_out = 8'h8D;
                    16'hB024: data_out = 8'h8C;
                    16'hB025: data_out = 8'h8B;
                    16'hB026: data_out = 8'h8A;
                    16'hB027: data_out = 8'h89;
                    16'hB028: data_out = 8'h88;
                    16'hB029: data_out = 8'h87;
                    16'hB02A: data_out = 8'h86;
                    16'hB02B: data_out = 8'h85;
                    16'hB02C: data_out = 8'h84;
                    16'hB02D: data_out = 8'h83;
                    16'hB02E: data_out = 8'h82;
                    16'hB02F: data_out = 8'h81;
                    16'hB030: data_out = 8'h0;
                    16'hB031: data_out = 8'h1;
                    16'hB032: data_out = 8'h2;
                    16'hB033: data_out = 8'h3;
                    16'hB034: data_out = 8'h4;
                    16'hB035: data_out = 8'h5;
                    16'hB036: data_out = 8'h6;
                    16'hB037: data_out = 8'h7;
                    16'hB038: data_out = 8'h8;
                    16'hB039: data_out = 8'h9;
                    16'hB03A: data_out = 8'hA;
                    16'hB03B: data_out = 8'hB;
                    16'hB03C: data_out = 8'hC;
                    16'hB03D: data_out = 8'hD;
                    16'hB03E: data_out = 8'hE;
                    16'hB03F: data_out = 8'hF;
                    16'hB040: data_out = 8'h10;
                    16'hB041: data_out = 8'h11;
                    16'hB042: data_out = 8'h12;
                    16'hB043: data_out = 8'h13;
                    16'hB044: data_out = 8'h14;
                    16'hB045: data_out = 8'h15;
                    16'hB046: data_out = 8'h16;
                    16'hB047: data_out = 8'h17;
                    16'hB048: data_out = 8'h18;
                    16'hB049: data_out = 8'h19;
                    16'hB04A: data_out = 8'h1A;
                    16'hB04B: data_out = 8'h1B;
                    16'hB04C: data_out = 8'h1C;
                    16'hB04D: data_out = 8'h1D;
                    16'hB04E: data_out = 8'h1E;
                    16'hB04F: data_out = 8'h1F;
                    16'hB050: data_out = 8'h20;
                    16'hB051: data_out = 8'h21;
                    16'hB052: data_out = 8'h22;
                    16'hB053: data_out = 8'h23;
                    16'hB054: data_out = 8'h24;
                    16'hB055: data_out = 8'h25;
                    16'hB056: data_out = 8'h26;
                    16'hB057: data_out = 8'h27;
                    16'hB058: data_out = 8'h28;
                    16'hB059: data_out = 8'h29;
                    16'hB05A: data_out = 8'h2A;
                    16'hB05B: data_out = 8'h2B;
                    16'hB05C: data_out = 8'h2C;
                    16'hB05D: data_out = 8'h2D;
                    16'hB05E: data_out = 8'h2E;
                    16'hB05F: data_out = 8'h2F;
                    16'hB060: data_out = 8'h30;
                    16'hB061: data_out = 8'h31;
                    16'hB062: data_out = 8'h32;
                    16'hB063: data_out = 8'h33;
                    16'hB064: data_out = 8'h34;
                    16'hB065: data_out = 8'h35;
                    16'hB066: data_out = 8'h36;
                    16'hB067: data_out = 8'h37;
                    16'hB068: data_out = 8'h38;
                    16'hB069: data_out = 8'h39;
                    16'hB06A: data_out = 8'h3A;
                    16'hB06B: data_out = 8'h3B;
                    16'hB06C: data_out = 8'h3C;
                    16'hB06D: data_out = 8'h3D;
                    16'hB06E: data_out = 8'h3E;
                    16'hB06F: data_out = 8'h3F;
                    16'hB070: data_out = 8'h40;
                    16'hB071: data_out = 8'h41;
                    16'hB072: data_out = 8'h42;
                    16'hB073: data_out = 8'h43;
                    16'hB074: data_out = 8'h44;
                    16'hB075: data_out = 8'h45;
                    16'hB076: data_out = 8'h46;
                    16'hB077: data_out = 8'h47;
                    16'hB078: data_out = 8'h48;
                    16'hB079: data_out = 8'h49;
                    16'hB07A: data_out = 8'h4A;
                    16'hB07B: data_out = 8'h4B;
                    16'hB07C: data_out = 8'h4C;
                    16'hB07D: data_out = 8'h4D;
                    16'hB07E: data_out = 8'h4E;
                    16'hB07F: data_out = 8'h4F;
                    16'hB080: data_out = 8'hB0;
                    16'hB081: data_out = 8'hB1;
                    16'hB082: data_out = 8'hB2;
                    16'hB083: data_out = 8'hB3;
                    16'hB084: data_out = 8'hB4;
                    16'hB085: data_out = 8'hB5;
                    16'hB086: data_out = 8'hB6;
                    16'hB087: data_out = 8'hB7;
                    16'hB088: data_out = 8'hB8;
                    16'hB089: data_out = 8'hB9;
                    16'hB08A: data_out = 8'hBA;
                    16'hB08B: data_out = 8'hBB;
                    16'hB08C: data_out = 8'hBC;
                    16'hB08D: data_out = 8'hBD;
                    16'hB08E: data_out = 8'hBE;
                    16'hB08F: data_out = 8'hBF;
                    16'hB090: data_out = 8'hC0;
                    16'hB091: data_out = 8'hC1;
                    16'hB092: data_out = 8'hC2;
                    16'hB093: data_out = 8'hC3;
                    16'hB094: data_out = 8'hC4;
                    16'hB095: data_out = 8'hC5;
                    16'hB096: data_out = 8'hC6;
                    16'hB097: data_out = 8'hC7;
                    16'hB098: data_out = 8'hC8;
                    16'hB099: data_out = 8'hC9;
                    16'hB09A: data_out = 8'hCA;
                    16'hB09B: data_out = 8'hCB;
                    16'hB09C: data_out = 8'hCC;
                    16'hB09D: data_out = 8'hCD;
                    16'hB09E: data_out = 8'hCE;
                    16'hB09F: data_out = 8'hCF;
                    16'hB0A0: data_out = 8'hD0;
                    16'hB0A1: data_out = 8'hD1;
                    16'hB0A2: data_out = 8'hD2;
                    16'hB0A3: data_out = 8'hD3;
                    16'hB0A4: data_out = 8'hD4;
                    16'hB0A5: data_out = 8'hD5;
                    16'hB0A6: data_out = 8'hD6;
                    16'hB0A7: data_out = 8'hD7;
                    16'hB0A8: data_out = 8'hD8;
                    16'hB0A9: data_out = 8'hD9;
                    16'hB0AA: data_out = 8'hDA;
                    16'hB0AB: data_out = 8'hDB;
                    16'hB0AC: data_out = 8'hDC;
                    16'hB0AD: data_out = 8'hDD;
                    16'hB0AE: data_out = 8'hDE;
                    16'hB0AF: data_out = 8'hDF;
                    16'hB0B0: data_out = 8'hE0;
                    16'hB0B1: data_out = 8'hE1;
                    16'hB0B2: data_out = 8'hE2;
                    16'hB0B3: data_out = 8'hE3;
                    16'hB0B4: data_out = 8'hE4;
                    16'hB0B5: data_out = 8'hE5;
                    16'hB0B6: data_out = 8'hE6;
                    16'hB0B7: data_out = 8'hE7;
                    16'hB0B8: data_out = 8'hE8;
                    16'hB0B9: data_out = 8'hE9;
                    16'hB0BA: data_out = 8'hEA;
                    16'hB0BB: data_out = 8'hEB;
                    16'hB0BC: data_out = 8'hEC;
                    16'hB0BD: data_out = 8'hED;
                    16'hB0BE: data_out = 8'hEE;
                    16'hB0BF: data_out = 8'hEF;
                    16'hB0C0: data_out = 8'hF0;
                    16'hB0C1: data_out = 8'hF1;
                    16'hB0C2: data_out = 8'hF2;
                    16'hB0C3: data_out = 8'hF3;
                    16'hB0C4: data_out = 8'hF4;
                    16'hB0C5: data_out = 8'hF5;
                    16'hB0C6: data_out = 8'hF6;
                    16'hB0C7: data_out = 8'hF7;
                    16'hB0C8: data_out = 8'hF8;
                    16'hB0C9: data_out = 8'hF9;
                    16'hB0CA: data_out = 8'hFA;
                    16'hB0CB: data_out = 8'hFB;
                    16'hB0CC: data_out = 8'hFC;
                    16'hB0CD: data_out = 8'hFD;
                    16'hB0CE: data_out = 8'hFE;
                    16'hB0CF: data_out = 8'hFF;
                    16'hB0D0: data_out = 8'h80;
                    16'hB0D1: data_out = 8'h81;
                    16'hB0D2: data_out = 8'h82;
                    16'hB0D3: data_out = 8'h83;
                    16'hB0D4: data_out = 8'h84;
                    16'hB0D5: data_out = 8'h85;
                    16'hB0D6: data_out = 8'h86;
                    16'hB0D7: data_out = 8'h87;
                    16'hB0D8: data_out = 8'h88;
                    16'hB0D9: data_out = 8'h89;
                    16'hB0DA: data_out = 8'h8A;
                    16'hB0DB: data_out = 8'h8B;
                    16'hB0DC: data_out = 8'h8C;
                    16'hB0DD: data_out = 8'h8D;
                    16'hB0DE: data_out = 8'h8E;
                    16'hB0DF: data_out = 8'h8F;
                    16'hB0E0: data_out = 8'h90;
                    16'hB0E1: data_out = 8'h91;
                    16'hB0E2: data_out = 8'h92;
                    16'hB0E3: data_out = 8'h93;
                    16'hB0E4: data_out = 8'h94;
                    16'hB0E5: data_out = 8'h95;
                    16'hB0E6: data_out = 8'h96;
                    16'hB0E7: data_out = 8'h97;
                    16'hB0E8: data_out = 8'h98;
                    16'hB0E9: data_out = 8'h99;
                    16'hB0EA: data_out = 8'h9A;
                    16'hB0EB: data_out = 8'h9B;
                    16'hB0EC: data_out = 8'h9C;
                    16'hB0ED: data_out = 8'h9D;
                    16'hB0EE: data_out = 8'h9E;
                    16'hB0EF: data_out = 8'h9F;
                    16'hB0F0: data_out = 8'hA0;
                    16'hB0F1: data_out = 8'hA1;
                    16'hB0F2: data_out = 8'hA2;
                    16'hB0F3: data_out = 8'hA3;
                    16'hB0F4: data_out = 8'hA4;
                    16'hB0F5: data_out = 8'hA5;
                    16'hB0F6: data_out = 8'hA6;
                    16'hB0F7: data_out = 8'hA7;
                    16'hB0F8: data_out = 8'hA8;
                    16'hB0F9: data_out = 8'hA9;
                    16'hB0FA: data_out = 8'hAA;
                    16'hB0FB: data_out = 8'hAB;
                    16'hB0FC: data_out = 8'hAC;
                    16'hB0FD: data_out = 8'hAD;
                    16'hB0FE: data_out = 8'hAE;
                    16'hB0FF: data_out = 8'hAF;
                    16'hB100: data_out = 8'hB1;
                    16'hB101: data_out = 8'hB0;
                    16'hB102: data_out = 8'hAF;
                    16'hB103: data_out = 8'hAE;
                    16'hB104: data_out = 8'hAD;
                    16'hB105: data_out = 8'hAC;
                    16'hB106: data_out = 8'hAB;
                    16'hB107: data_out = 8'hAA;
                    16'hB108: data_out = 8'hA9;
                    16'hB109: data_out = 8'hA8;
                    16'hB10A: data_out = 8'hA7;
                    16'hB10B: data_out = 8'hA6;
                    16'hB10C: data_out = 8'hA5;
                    16'hB10D: data_out = 8'hA4;
                    16'hB10E: data_out = 8'hA3;
                    16'hB10F: data_out = 8'hA2;
                    16'hB110: data_out = 8'hA1;
                    16'hB111: data_out = 8'hA0;
                    16'hB112: data_out = 8'h9F;
                    16'hB113: data_out = 8'h9E;
                    16'hB114: data_out = 8'h9D;
                    16'hB115: data_out = 8'h9C;
                    16'hB116: data_out = 8'h9B;
                    16'hB117: data_out = 8'h9A;
                    16'hB118: data_out = 8'h99;
                    16'hB119: data_out = 8'h98;
                    16'hB11A: data_out = 8'h97;
                    16'hB11B: data_out = 8'h96;
                    16'hB11C: data_out = 8'h95;
                    16'hB11D: data_out = 8'h94;
                    16'hB11E: data_out = 8'h93;
                    16'hB11F: data_out = 8'h92;
                    16'hB120: data_out = 8'h91;
                    16'hB121: data_out = 8'h90;
                    16'hB122: data_out = 8'h8F;
                    16'hB123: data_out = 8'h8E;
                    16'hB124: data_out = 8'h8D;
                    16'hB125: data_out = 8'h8C;
                    16'hB126: data_out = 8'h8B;
                    16'hB127: data_out = 8'h8A;
                    16'hB128: data_out = 8'h89;
                    16'hB129: data_out = 8'h88;
                    16'hB12A: data_out = 8'h87;
                    16'hB12B: data_out = 8'h86;
                    16'hB12C: data_out = 8'h85;
                    16'hB12D: data_out = 8'h84;
                    16'hB12E: data_out = 8'h83;
                    16'hB12F: data_out = 8'h82;
                    16'hB130: data_out = 8'h81;
                    16'hB131: data_out = 8'h0;
                    16'hB132: data_out = 8'h1;
                    16'hB133: data_out = 8'h2;
                    16'hB134: data_out = 8'h3;
                    16'hB135: data_out = 8'h4;
                    16'hB136: data_out = 8'h5;
                    16'hB137: data_out = 8'h6;
                    16'hB138: data_out = 8'h7;
                    16'hB139: data_out = 8'h8;
                    16'hB13A: data_out = 8'h9;
                    16'hB13B: data_out = 8'hA;
                    16'hB13C: data_out = 8'hB;
                    16'hB13D: data_out = 8'hC;
                    16'hB13E: data_out = 8'hD;
                    16'hB13F: data_out = 8'hE;
                    16'hB140: data_out = 8'hF;
                    16'hB141: data_out = 8'h10;
                    16'hB142: data_out = 8'h11;
                    16'hB143: data_out = 8'h12;
                    16'hB144: data_out = 8'h13;
                    16'hB145: data_out = 8'h14;
                    16'hB146: data_out = 8'h15;
                    16'hB147: data_out = 8'h16;
                    16'hB148: data_out = 8'h17;
                    16'hB149: data_out = 8'h18;
                    16'hB14A: data_out = 8'h19;
                    16'hB14B: data_out = 8'h1A;
                    16'hB14C: data_out = 8'h1B;
                    16'hB14D: data_out = 8'h1C;
                    16'hB14E: data_out = 8'h1D;
                    16'hB14F: data_out = 8'h1E;
                    16'hB150: data_out = 8'h1F;
                    16'hB151: data_out = 8'h20;
                    16'hB152: data_out = 8'h21;
                    16'hB153: data_out = 8'h22;
                    16'hB154: data_out = 8'h23;
                    16'hB155: data_out = 8'h24;
                    16'hB156: data_out = 8'h25;
                    16'hB157: data_out = 8'h26;
                    16'hB158: data_out = 8'h27;
                    16'hB159: data_out = 8'h28;
                    16'hB15A: data_out = 8'h29;
                    16'hB15B: data_out = 8'h2A;
                    16'hB15C: data_out = 8'h2B;
                    16'hB15D: data_out = 8'h2C;
                    16'hB15E: data_out = 8'h2D;
                    16'hB15F: data_out = 8'h2E;
                    16'hB160: data_out = 8'h2F;
                    16'hB161: data_out = 8'h30;
                    16'hB162: data_out = 8'h31;
                    16'hB163: data_out = 8'h32;
                    16'hB164: data_out = 8'h33;
                    16'hB165: data_out = 8'h34;
                    16'hB166: data_out = 8'h35;
                    16'hB167: data_out = 8'h36;
                    16'hB168: data_out = 8'h37;
                    16'hB169: data_out = 8'h38;
                    16'hB16A: data_out = 8'h39;
                    16'hB16B: data_out = 8'h3A;
                    16'hB16C: data_out = 8'h3B;
                    16'hB16D: data_out = 8'h3C;
                    16'hB16E: data_out = 8'h3D;
                    16'hB16F: data_out = 8'h3E;
                    16'hB170: data_out = 8'h3F;
                    16'hB171: data_out = 8'h40;
                    16'hB172: data_out = 8'h41;
                    16'hB173: data_out = 8'h42;
                    16'hB174: data_out = 8'h43;
                    16'hB175: data_out = 8'h44;
                    16'hB176: data_out = 8'h45;
                    16'hB177: data_out = 8'h46;
                    16'hB178: data_out = 8'h47;
                    16'hB179: data_out = 8'h48;
                    16'hB17A: data_out = 8'h49;
                    16'hB17B: data_out = 8'h4A;
                    16'hB17C: data_out = 8'h4B;
                    16'hB17D: data_out = 8'h4C;
                    16'hB17E: data_out = 8'h4D;
                    16'hB17F: data_out = 8'h4E;
                    16'hB180: data_out = 8'hB1;
                    16'hB181: data_out = 8'hB2;
                    16'hB182: data_out = 8'hB3;
                    16'hB183: data_out = 8'hB4;
                    16'hB184: data_out = 8'hB5;
                    16'hB185: data_out = 8'hB6;
                    16'hB186: data_out = 8'hB7;
                    16'hB187: data_out = 8'hB8;
                    16'hB188: data_out = 8'hB9;
                    16'hB189: data_out = 8'hBA;
                    16'hB18A: data_out = 8'hBB;
                    16'hB18B: data_out = 8'hBC;
                    16'hB18C: data_out = 8'hBD;
                    16'hB18D: data_out = 8'hBE;
                    16'hB18E: data_out = 8'hBF;
                    16'hB18F: data_out = 8'hC0;
                    16'hB190: data_out = 8'hC1;
                    16'hB191: data_out = 8'hC2;
                    16'hB192: data_out = 8'hC3;
                    16'hB193: data_out = 8'hC4;
                    16'hB194: data_out = 8'hC5;
                    16'hB195: data_out = 8'hC6;
                    16'hB196: data_out = 8'hC7;
                    16'hB197: data_out = 8'hC8;
                    16'hB198: data_out = 8'hC9;
                    16'hB199: data_out = 8'hCA;
                    16'hB19A: data_out = 8'hCB;
                    16'hB19B: data_out = 8'hCC;
                    16'hB19C: data_out = 8'hCD;
                    16'hB19D: data_out = 8'hCE;
                    16'hB19E: data_out = 8'hCF;
                    16'hB19F: data_out = 8'hD0;
                    16'hB1A0: data_out = 8'hD1;
                    16'hB1A1: data_out = 8'hD2;
                    16'hB1A2: data_out = 8'hD3;
                    16'hB1A3: data_out = 8'hD4;
                    16'hB1A4: data_out = 8'hD5;
                    16'hB1A5: data_out = 8'hD6;
                    16'hB1A6: data_out = 8'hD7;
                    16'hB1A7: data_out = 8'hD8;
                    16'hB1A8: data_out = 8'hD9;
                    16'hB1A9: data_out = 8'hDA;
                    16'hB1AA: data_out = 8'hDB;
                    16'hB1AB: data_out = 8'hDC;
                    16'hB1AC: data_out = 8'hDD;
                    16'hB1AD: data_out = 8'hDE;
                    16'hB1AE: data_out = 8'hDF;
                    16'hB1AF: data_out = 8'hE0;
                    16'hB1B0: data_out = 8'hE1;
                    16'hB1B1: data_out = 8'hE2;
                    16'hB1B2: data_out = 8'hE3;
                    16'hB1B3: data_out = 8'hE4;
                    16'hB1B4: data_out = 8'hE5;
                    16'hB1B5: data_out = 8'hE6;
                    16'hB1B6: data_out = 8'hE7;
                    16'hB1B7: data_out = 8'hE8;
                    16'hB1B8: data_out = 8'hE9;
                    16'hB1B9: data_out = 8'hEA;
                    16'hB1BA: data_out = 8'hEB;
                    16'hB1BB: data_out = 8'hEC;
                    16'hB1BC: data_out = 8'hED;
                    16'hB1BD: data_out = 8'hEE;
                    16'hB1BE: data_out = 8'hEF;
                    16'hB1BF: data_out = 8'hF0;
                    16'hB1C0: data_out = 8'hF1;
                    16'hB1C1: data_out = 8'hF2;
                    16'hB1C2: data_out = 8'hF3;
                    16'hB1C3: data_out = 8'hF4;
                    16'hB1C4: data_out = 8'hF5;
                    16'hB1C5: data_out = 8'hF6;
                    16'hB1C6: data_out = 8'hF7;
                    16'hB1C7: data_out = 8'hF8;
                    16'hB1C8: data_out = 8'hF9;
                    16'hB1C9: data_out = 8'hFA;
                    16'hB1CA: data_out = 8'hFB;
                    16'hB1CB: data_out = 8'hFC;
                    16'hB1CC: data_out = 8'hFD;
                    16'hB1CD: data_out = 8'hFE;
                    16'hB1CE: data_out = 8'hFF;
                    16'hB1CF: data_out = 8'h80;
                    16'hB1D0: data_out = 8'h81;
                    16'hB1D1: data_out = 8'h82;
                    16'hB1D2: data_out = 8'h83;
                    16'hB1D3: data_out = 8'h84;
                    16'hB1D4: data_out = 8'h85;
                    16'hB1D5: data_out = 8'h86;
                    16'hB1D6: data_out = 8'h87;
                    16'hB1D7: data_out = 8'h88;
                    16'hB1D8: data_out = 8'h89;
                    16'hB1D9: data_out = 8'h8A;
                    16'hB1DA: data_out = 8'h8B;
                    16'hB1DB: data_out = 8'h8C;
                    16'hB1DC: data_out = 8'h8D;
                    16'hB1DD: data_out = 8'h8E;
                    16'hB1DE: data_out = 8'h8F;
                    16'hB1DF: data_out = 8'h90;
                    16'hB1E0: data_out = 8'h91;
                    16'hB1E1: data_out = 8'h92;
                    16'hB1E2: data_out = 8'h93;
                    16'hB1E3: data_out = 8'h94;
                    16'hB1E4: data_out = 8'h95;
                    16'hB1E5: data_out = 8'h96;
                    16'hB1E6: data_out = 8'h97;
                    16'hB1E7: data_out = 8'h98;
                    16'hB1E8: data_out = 8'h99;
                    16'hB1E9: data_out = 8'h9A;
                    16'hB1EA: data_out = 8'h9B;
                    16'hB1EB: data_out = 8'h9C;
                    16'hB1EC: data_out = 8'h9D;
                    16'hB1ED: data_out = 8'h9E;
                    16'hB1EE: data_out = 8'h9F;
                    16'hB1EF: data_out = 8'hA0;
                    16'hB1F0: data_out = 8'hA1;
                    16'hB1F1: data_out = 8'hA2;
                    16'hB1F2: data_out = 8'hA3;
                    16'hB1F3: data_out = 8'hA4;
                    16'hB1F4: data_out = 8'hA5;
                    16'hB1F5: data_out = 8'hA6;
                    16'hB1F6: data_out = 8'hA7;
                    16'hB1F7: data_out = 8'hA8;
                    16'hB1F8: data_out = 8'hA9;
                    16'hB1F9: data_out = 8'hAA;
                    16'hB1FA: data_out = 8'hAB;
                    16'hB1FB: data_out = 8'hAC;
                    16'hB1FC: data_out = 8'hAD;
                    16'hB1FD: data_out = 8'hAE;
                    16'hB1FE: data_out = 8'hAF;
                    16'hB1FF: data_out = 8'hB0;
                    16'hB200: data_out = 8'hB2;
                    16'hB201: data_out = 8'hB1;
                    16'hB202: data_out = 8'hB0;
                    16'hB203: data_out = 8'hAF;
                    16'hB204: data_out = 8'hAE;
                    16'hB205: data_out = 8'hAD;
                    16'hB206: data_out = 8'hAC;
                    16'hB207: data_out = 8'hAB;
                    16'hB208: data_out = 8'hAA;
                    16'hB209: data_out = 8'hA9;
                    16'hB20A: data_out = 8'hA8;
                    16'hB20B: data_out = 8'hA7;
                    16'hB20C: data_out = 8'hA6;
                    16'hB20D: data_out = 8'hA5;
                    16'hB20E: data_out = 8'hA4;
                    16'hB20F: data_out = 8'hA3;
                    16'hB210: data_out = 8'hA2;
                    16'hB211: data_out = 8'hA1;
                    16'hB212: data_out = 8'hA0;
                    16'hB213: data_out = 8'h9F;
                    16'hB214: data_out = 8'h9E;
                    16'hB215: data_out = 8'h9D;
                    16'hB216: data_out = 8'h9C;
                    16'hB217: data_out = 8'h9B;
                    16'hB218: data_out = 8'h9A;
                    16'hB219: data_out = 8'h99;
                    16'hB21A: data_out = 8'h98;
                    16'hB21B: data_out = 8'h97;
                    16'hB21C: data_out = 8'h96;
                    16'hB21D: data_out = 8'h95;
                    16'hB21E: data_out = 8'h94;
                    16'hB21F: data_out = 8'h93;
                    16'hB220: data_out = 8'h92;
                    16'hB221: data_out = 8'h91;
                    16'hB222: data_out = 8'h90;
                    16'hB223: data_out = 8'h8F;
                    16'hB224: data_out = 8'h8E;
                    16'hB225: data_out = 8'h8D;
                    16'hB226: data_out = 8'h8C;
                    16'hB227: data_out = 8'h8B;
                    16'hB228: data_out = 8'h8A;
                    16'hB229: data_out = 8'h89;
                    16'hB22A: data_out = 8'h88;
                    16'hB22B: data_out = 8'h87;
                    16'hB22C: data_out = 8'h86;
                    16'hB22D: data_out = 8'h85;
                    16'hB22E: data_out = 8'h84;
                    16'hB22F: data_out = 8'h83;
                    16'hB230: data_out = 8'h82;
                    16'hB231: data_out = 8'h81;
                    16'hB232: data_out = 8'h0;
                    16'hB233: data_out = 8'h1;
                    16'hB234: data_out = 8'h2;
                    16'hB235: data_out = 8'h3;
                    16'hB236: data_out = 8'h4;
                    16'hB237: data_out = 8'h5;
                    16'hB238: data_out = 8'h6;
                    16'hB239: data_out = 8'h7;
                    16'hB23A: data_out = 8'h8;
                    16'hB23B: data_out = 8'h9;
                    16'hB23C: data_out = 8'hA;
                    16'hB23D: data_out = 8'hB;
                    16'hB23E: data_out = 8'hC;
                    16'hB23F: data_out = 8'hD;
                    16'hB240: data_out = 8'hE;
                    16'hB241: data_out = 8'hF;
                    16'hB242: data_out = 8'h10;
                    16'hB243: data_out = 8'h11;
                    16'hB244: data_out = 8'h12;
                    16'hB245: data_out = 8'h13;
                    16'hB246: data_out = 8'h14;
                    16'hB247: data_out = 8'h15;
                    16'hB248: data_out = 8'h16;
                    16'hB249: data_out = 8'h17;
                    16'hB24A: data_out = 8'h18;
                    16'hB24B: data_out = 8'h19;
                    16'hB24C: data_out = 8'h1A;
                    16'hB24D: data_out = 8'h1B;
                    16'hB24E: data_out = 8'h1C;
                    16'hB24F: data_out = 8'h1D;
                    16'hB250: data_out = 8'h1E;
                    16'hB251: data_out = 8'h1F;
                    16'hB252: data_out = 8'h20;
                    16'hB253: data_out = 8'h21;
                    16'hB254: data_out = 8'h22;
                    16'hB255: data_out = 8'h23;
                    16'hB256: data_out = 8'h24;
                    16'hB257: data_out = 8'h25;
                    16'hB258: data_out = 8'h26;
                    16'hB259: data_out = 8'h27;
                    16'hB25A: data_out = 8'h28;
                    16'hB25B: data_out = 8'h29;
                    16'hB25C: data_out = 8'h2A;
                    16'hB25D: data_out = 8'h2B;
                    16'hB25E: data_out = 8'h2C;
                    16'hB25F: data_out = 8'h2D;
                    16'hB260: data_out = 8'h2E;
                    16'hB261: data_out = 8'h2F;
                    16'hB262: data_out = 8'h30;
                    16'hB263: data_out = 8'h31;
                    16'hB264: data_out = 8'h32;
                    16'hB265: data_out = 8'h33;
                    16'hB266: data_out = 8'h34;
                    16'hB267: data_out = 8'h35;
                    16'hB268: data_out = 8'h36;
                    16'hB269: data_out = 8'h37;
                    16'hB26A: data_out = 8'h38;
                    16'hB26B: data_out = 8'h39;
                    16'hB26C: data_out = 8'h3A;
                    16'hB26D: data_out = 8'h3B;
                    16'hB26E: data_out = 8'h3C;
                    16'hB26F: data_out = 8'h3D;
                    16'hB270: data_out = 8'h3E;
                    16'hB271: data_out = 8'h3F;
                    16'hB272: data_out = 8'h40;
                    16'hB273: data_out = 8'h41;
                    16'hB274: data_out = 8'h42;
                    16'hB275: data_out = 8'h43;
                    16'hB276: data_out = 8'h44;
                    16'hB277: data_out = 8'h45;
                    16'hB278: data_out = 8'h46;
                    16'hB279: data_out = 8'h47;
                    16'hB27A: data_out = 8'h48;
                    16'hB27B: data_out = 8'h49;
                    16'hB27C: data_out = 8'h4A;
                    16'hB27D: data_out = 8'h4B;
                    16'hB27E: data_out = 8'h4C;
                    16'hB27F: data_out = 8'h4D;
                    16'hB280: data_out = 8'hB2;
                    16'hB281: data_out = 8'hB3;
                    16'hB282: data_out = 8'hB4;
                    16'hB283: data_out = 8'hB5;
                    16'hB284: data_out = 8'hB6;
                    16'hB285: data_out = 8'hB7;
                    16'hB286: data_out = 8'hB8;
                    16'hB287: data_out = 8'hB9;
                    16'hB288: data_out = 8'hBA;
                    16'hB289: data_out = 8'hBB;
                    16'hB28A: data_out = 8'hBC;
                    16'hB28B: data_out = 8'hBD;
                    16'hB28C: data_out = 8'hBE;
                    16'hB28D: data_out = 8'hBF;
                    16'hB28E: data_out = 8'hC0;
                    16'hB28F: data_out = 8'hC1;
                    16'hB290: data_out = 8'hC2;
                    16'hB291: data_out = 8'hC3;
                    16'hB292: data_out = 8'hC4;
                    16'hB293: data_out = 8'hC5;
                    16'hB294: data_out = 8'hC6;
                    16'hB295: data_out = 8'hC7;
                    16'hB296: data_out = 8'hC8;
                    16'hB297: data_out = 8'hC9;
                    16'hB298: data_out = 8'hCA;
                    16'hB299: data_out = 8'hCB;
                    16'hB29A: data_out = 8'hCC;
                    16'hB29B: data_out = 8'hCD;
                    16'hB29C: data_out = 8'hCE;
                    16'hB29D: data_out = 8'hCF;
                    16'hB29E: data_out = 8'hD0;
                    16'hB29F: data_out = 8'hD1;
                    16'hB2A0: data_out = 8'hD2;
                    16'hB2A1: data_out = 8'hD3;
                    16'hB2A2: data_out = 8'hD4;
                    16'hB2A3: data_out = 8'hD5;
                    16'hB2A4: data_out = 8'hD6;
                    16'hB2A5: data_out = 8'hD7;
                    16'hB2A6: data_out = 8'hD8;
                    16'hB2A7: data_out = 8'hD9;
                    16'hB2A8: data_out = 8'hDA;
                    16'hB2A9: data_out = 8'hDB;
                    16'hB2AA: data_out = 8'hDC;
                    16'hB2AB: data_out = 8'hDD;
                    16'hB2AC: data_out = 8'hDE;
                    16'hB2AD: data_out = 8'hDF;
                    16'hB2AE: data_out = 8'hE0;
                    16'hB2AF: data_out = 8'hE1;
                    16'hB2B0: data_out = 8'hE2;
                    16'hB2B1: data_out = 8'hE3;
                    16'hB2B2: data_out = 8'hE4;
                    16'hB2B3: data_out = 8'hE5;
                    16'hB2B4: data_out = 8'hE6;
                    16'hB2B5: data_out = 8'hE7;
                    16'hB2B6: data_out = 8'hE8;
                    16'hB2B7: data_out = 8'hE9;
                    16'hB2B8: data_out = 8'hEA;
                    16'hB2B9: data_out = 8'hEB;
                    16'hB2BA: data_out = 8'hEC;
                    16'hB2BB: data_out = 8'hED;
                    16'hB2BC: data_out = 8'hEE;
                    16'hB2BD: data_out = 8'hEF;
                    16'hB2BE: data_out = 8'hF0;
                    16'hB2BF: data_out = 8'hF1;
                    16'hB2C0: data_out = 8'hF2;
                    16'hB2C1: data_out = 8'hF3;
                    16'hB2C2: data_out = 8'hF4;
                    16'hB2C3: data_out = 8'hF5;
                    16'hB2C4: data_out = 8'hF6;
                    16'hB2C5: data_out = 8'hF7;
                    16'hB2C6: data_out = 8'hF8;
                    16'hB2C7: data_out = 8'hF9;
                    16'hB2C8: data_out = 8'hFA;
                    16'hB2C9: data_out = 8'hFB;
                    16'hB2CA: data_out = 8'hFC;
                    16'hB2CB: data_out = 8'hFD;
                    16'hB2CC: data_out = 8'hFE;
                    16'hB2CD: data_out = 8'hFF;
                    16'hB2CE: data_out = 8'h80;
                    16'hB2CF: data_out = 8'h81;
                    16'hB2D0: data_out = 8'h82;
                    16'hB2D1: data_out = 8'h83;
                    16'hB2D2: data_out = 8'h84;
                    16'hB2D3: data_out = 8'h85;
                    16'hB2D4: data_out = 8'h86;
                    16'hB2D5: data_out = 8'h87;
                    16'hB2D6: data_out = 8'h88;
                    16'hB2D7: data_out = 8'h89;
                    16'hB2D8: data_out = 8'h8A;
                    16'hB2D9: data_out = 8'h8B;
                    16'hB2DA: data_out = 8'h8C;
                    16'hB2DB: data_out = 8'h8D;
                    16'hB2DC: data_out = 8'h8E;
                    16'hB2DD: data_out = 8'h8F;
                    16'hB2DE: data_out = 8'h90;
                    16'hB2DF: data_out = 8'h91;
                    16'hB2E0: data_out = 8'h92;
                    16'hB2E1: data_out = 8'h93;
                    16'hB2E2: data_out = 8'h94;
                    16'hB2E3: data_out = 8'h95;
                    16'hB2E4: data_out = 8'h96;
                    16'hB2E5: data_out = 8'h97;
                    16'hB2E6: data_out = 8'h98;
                    16'hB2E7: data_out = 8'h99;
                    16'hB2E8: data_out = 8'h9A;
                    16'hB2E9: data_out = 8'h9B;
                    16'hB2EA: data_out = 8'h9C;
                    16'hB2EB: data_out = 8'h9D;
                    16'hB2EC: data_out = 8'h9E;
                    16'hB2ED: data_out = 8'h9F;
                    16'hB2EE: data_out = 8'hA0;
                    16'hB2EF: data_out = 8'hA1;
                    16'hB2F0: data_out = 8'hA2;
                    16'hB2F1: data_out = 8'hA3;
                    16'hB2F2: data_out = 8'hA4;
                    16'hB2F3: data_out = 8'hA5;
                    16'hB2F4: data_out = 8'hA6;
                    16'hB2F5: data_out = 8'hA7;
                    16'hB2F6: data_out = 8'hA8;
                    16'hB2F7: data_out = 8'hA9;
                    16'hB2F8: data_out = 8'hAA;
                    16'hB2F9: data_out = 8'hAB;
                    16'hB2FA: data_out = 8'hAC;
                    16'hB2FB: data_out = 8'hAD;
                    16'hB2FC: data_out = 8'hAE;
                    16'hB2FD: data_out = 8'hAF;
                    16'hB2FE: data_out = 8'hB0;
                    16'hB2FF: data_out = 8'hB1;
                    16'hB300: data_out = 8'hB3;
                    16'hB301: data_out = 8'hB2;
                    16'hB302: data_out = 8'hB1;
                    16'hB303: data_out = 8'hB0;
                    16'hB304: data_out = 8'hAF;
                    16'hB305: data_out = 8'hAE;
                    16'hB306: data_out = 8'hAD;
                    16'hB307: data_out = 8'hAC;
                    16'hB308: data_out = 8'hAB;
                    16'hB309: data_out = 8'hAA;
                    16'hB30A: data_out = 8'hA9;
                    16'hB30B: data_out = 8'hA8;
                    16'hB30C: data_out = 8'hA7;
                    16'hB30D: data_out = 8'hA6;
                    16'hB30E: data_out = 8'hA5;
                    16'hB30F: data_out = 8'hA4;
                    16'hB310: data_out = 8'hA3;
                    16'hB311: data_out = 8'hA2;
                    16'hB312: data_out = 8'hA1;
                    16'hB313: data_out = 8'hA0;
                    16'hB314: data_out = 8'h9F;
                    16'hB315: data_out = 8'h9E;
                    16'hB316: data_out = 8'h9D;
                    16'hB317: data_out = 8'h9C;
                    16'hB318: data_out = 8'h9B;
                    16'hB319: data_out = 8'h9A;
                    16'hB31A: data_out = 8'h99;
                    16'hB31B: data_out = 8'h98;
                    16'hB31C: data_out = 8'h97;
                    16'hB31D: data_out = 8'h96;
                    16'hB31E: data_out = 8'h95;
                    16'hB31F: data_out = 8'h94;
                    16'hB320: data_out = 8'h93;
                    16'hB321: data_out = 8'h92;
                    16'hB322: data_out = 8'h91;
                    16'hB323: data_out = 8'h90;
                    16'hB324: data_out = 8'h8F;
                    16'hB325: data_out = 8'h8E;
                    16'hB326: data_out = 8'h8D;
                    16'hB327: data_out = 8'h8C;
                    16'hB328: data_out = 8'h8B;
                    16'hB329: data_out = 8'h8A;
                    16'hB32A: data_out = 8'h89;
                    16'hB32B: data_out = 8'h88;
                    16'hB32C: data_out = 8'h87;
                    16'hB32D: data_out = 8'h86;
                    16'hB32E: data_out = 8'h85;
                    16'hB32F: data_out = 8'h84;
                    16'hB330: data_out = 8'h83;
                    16'hB331: data_out = 8'h82;
                    16'hB332: data_out = 8'h81;
                    16'hB333: data_out = 8'h0;
                    16'hB334: data_out = 8'h1;
                    16'hB335: data_out = 8'h2;
                    16'hB336: data_out = 8'h3;
                    16'hB337: data_out = 8'h4;
                    16'hB338: data_out = 8'h5;
                    16'hB339: data_out = 8'h6;
                    16'hB33A: data_out = 8'h7;
                    16'hB33B: data_out = 8'h8;
                    16'hB33C: data_out = 8'h9;
                    16'hB33D: data_out = 8'hA;
                    16'hB33E: data_out = 8'hB;
                    16'hB33F: data_out = 8'hC;
                    16'hB340: data_out = 8'hD;
                    16'hB341: data_out = 8'hE;
                    16'hB342: data_out = 8'hF;
                    16'hB343: data_out = 8'h10;
                    16'hB344: data_out = 8'h11;
                    16'hB345: data_out = 8'h12;
                    16'hB346: data_out = 8'h13;
                    16'hB347: data_out = 8'h14;
                    16'hB348: data_out = 8'h15;
                    16'hB349: data_out = 8'h16;
                    16'hB34A: data_out = 8'h17;
                    16'hB34B: data_out = 8'h18;
                    16'hB34C: data_out = 8'h19;
                    16'hB34D: data_out = 8'h1A;
                    16'hB34E: data_out = 8'h1B;
                    16'hB34F: data_out = 8'h1C;
                    16'hB350: data_out = 8'h1D;
                    16'hB351: data_out = 8'h1E;
                    16'hB352: data_out = 8'h1F;
                    16'hB353: data_out = 8'h20;
                    16'hB354: data_out = 8'h21;
                    16'hB355: data_out = 8'h22;
                    16'hB356: data_out = 8'h23;
                    16'hB357: data_out = 8'h24;
                    16'hB358: data_out = 8'h25;
                    16'hB359: data_out = 8'h26;
                    16'hB35A: data_out = 8'h27;
                    16'hB35B: data_out = 8'h28;
                    16'hB35C: data_out = 8'h29;
                    16'hB35D: data_out = 8'h2A;
                    16'hB35E: data_out = 8'h2B;
                    16'hB35F: data_out = 8'h2C;
                    16'hB360: data_out = 8'h2D;
                    16'hB361: data_out = 8'h2E;
                    16'hB362: data_out = 8'h2F;
                    16'hB363: data_out = 8'h30;
                    16'hB364: data_out = 8'h31;
                    16'hB365: data_out = 8'h32;
                    16'hB366: data_out = 8'h33;
                    16'hB367: data_out = 8'h34;
                    16'hB368: data_out = 8'h35;
                    16'hB369: data_out = 8'h36;
                    16'hB36A: data_out = 8'h37;
                    16'hB36B: data_out = 8'h38;
                    16'hB36C: data_out = 8'h39;
                    16'hB36D: data_out = 8'h3A;
                    16'hB36E: data_out = 8'h3B;
                    16'hB36F: data_out = 8'h3C;
                    16'hB370: data_out = 8'h3D;
                    16'hB371: data_out = 8'h3E;
                    16'hB372: data_out = 8'h3F;
                    16'hB373: data_out = 8'h40;
                    16'hB374: data_out = 8'h41;
                    16'hB375: data_out = 8'h42;
                    16'hB376: data_out = 8'h43;
                    16'hB377: data_out = 8'h44;
                    16'hB378: data_out = 8'h45;
                    16'hB379: data_out = 8'h46;
                    16'hB37A: data_out = 8'h47;
                    16'hB37B: data_out = 8'h48;
                    16'hB37C: data_out = 8'h49;
                    16'hB37D: data_out = 8'h4A;
                    16'hB37E: data_out = 8'h4B;
                    16'hB37F: data_out = 8'h4C;
                    16'hB380: data_out = 8'hB3;
                    16'hB381: data_out = 8'hB4;
                    16'hB382: data_out = 8'hB5;
                    16'hB383: data_out = 8'hB6;
                    16'hB384: data_out = 8'hB7;
                    16'hB385: data_out = 8'hB8;
                    16'hB386: data_out = 8'hB9;
                    16'hB387: data_out = 8'hBA;
                    16'hB388: data_out = 8'hBB;
                    16'hB389: data_out = 8'hBC;
                    16'hB38A: data_out = 8'hBD;
                    16'hB38B: data_out = 8'hBE;
                    16'hB38C: data_out = 8'hBF;
                    16'hB38D: data_out = 8'hC0;
                    16'hB38E: data_out = 8'hC1;
                    16'hB38F: data_out = 8'hC2;
                    16'hB390: data_out = 8'hC3;
                    16'hB391: data_out = 8'hC4;
                    16'hB392: data_out = 8'hC5;
                    16'hB393: data_out = 8'hC6;
                    16'hB394: data_out = 8'hC7;
                    16'hB395: data_out = 8'hC8;
                    16'hB396: data_out = 8'hC9;
                    16'hB397: data_out = 8'hCA;
                    16'hB398: data_out = 8'hCB;
                    16'hB399: data_out = 8'hCC;
                    16'hB39A: data_out = 8'hCD;
                    16'hB39B: data_out = 8'hCE;
                    16'hB39C: data_out = 8'hCF;
                    16'hB39D: data_out = 8'hD0;
                    16'hB39E: data_out = 8'hD1;
                    16'hB39F: data_out = 8'hD2;
                    16'hB3A0: data_out = 8'hD3;
                    16'hB3A1: data_out = 8'hD4;
                    16'hB3A2: data_out = 8'hD5;
                    16'hB3A3: data_out = 8'hD6;
                    16'hB3A4: data_out = 8'hD7;
                    16'hB3A5: data_out = 8'hD8;
                    16'hB3A6: data_out = 8'hD9;
                    16'hB3A7: data_out = 8'hDA;
                    16'hB3A8: data_out = 8'hDB;
                    16'hB3A9: data_out = 8'hDC;
                    16'hB3AA: data_out = 8'hDD;
                    16'hB3AB: data_out = 8'hDE;
                    16'hB3AC: data_out = 8'hDF;
                    16'hB3AD: data_out = 8'hE0;
                    16'hB3AE: data_out = 8'hE1;
                    16'hB3AF: data_out = 8'hE2;
                    16'hB3B0: data_out = 8'hE3;
                    16'hB3B1: data_out = 8'hE4;
                    16'hB3B2: data_out = 8'hE5;
                    16'hB3B3: data_out = 8'hE6;
                    16'hB3B4: data_out = 8'hE7;
                    16'hB3B5: data_out = 8'hE8;
                    16'hB3B6: data_out = 8'hE9;
                    16'hB3B7: data_out = 8'hEA;
                    16'hB3B8: data_out = 8'hEB;
                    16'hB3B9: data_out = 8'hEC;
                    16'hB3BA: data_out = 8'hED;
                    16'hB3BB: data_out = 8'hEE;
                    16'hB3BC: data_out = 8'hEF;
                    16'hB3BD: data_out = 8'hF0;
                    16'hB3BE: data_out = 8'hF1;
                    16'hB3BF: data_out = 8'hF2;
                    16'hB3C0: data_out = 8'hF3;
                    16'hB3C1: data_out = 8'hF4;
                    16'hB3C2: data_out = 8'hF5;
                    16'hB3C3: data_out = 8'hF6;
                    16'hB3C4: data_out = 8'hF7;
                    16'hB3C5: data_out = 8'hF8;
                    16'hB3C6: data_out = 8'hF9;
                    16'hB3C7: data_out = 8'hFA;
                    16'hB3C8: data_out = 8'hFB;
                    16'hB3C9: data_out = 8'hFC;
                    16'hB3CA: data_out = 8'hFD;
                    16'hB3CB: data_out = 8'hFE;
                    16'hB3CC: data_out = 8'hFF;
                    16'hB3CD: data_out = 8'h80;
                    16'hB3CE: data_out = 8'h81;
                    16'hB3CF: data_out = 8'h82;
                    16'hB3D0: data_out = 8'h83;
                    16'hB3D1: data_out = 8'h84;
                    16'hB3D2: data_out = 8'h85;
                    16'hB3D3: data_out = 8'h86;
                    16'hB3D4: data_out = 8'h87;
                    16'hB3D5: data_out = 8'h88;
                    16'hB3D6: data_out = 8'h89;
                    16'hB3D7: data_out = 8'h8A;
                    16'hB3D8: data_out = 8'h8B;
                    16'hB3D9: data_out = 8'h8C;
                    16'hB3DA: data_out = 8'h8D;
                    16'hB3DB: data_out = 8'h8E;
                    16'hB3DC: data_out = 8'h8F;
                    16'hB3DD: data_out = 8'h90;
                    16'hB3DE: data_out = 8'h91;
                    16'hB3DF: data_out = 8'h92;
                    16'hB3E0: data_out = 8'h93;
                    16'hB3E1: data_out = 8'h94;
                    16'hB3E2: data_out = 8'h95;
                    16'hB3E3: data_out = 8'h96;
                    16'hB3E4: data_out = 8'h97;
                    16'hB3E5: data_out = 8'h98;
                    16'hB3E6: data_out = 8'h99;
                    16'hB3E7: data_out = 8'h9A;
                    16'hB3E8: data_out = 8'h9B;
                    16'hB3E9: data_out = 8'h9C;
                    16'hB3EA: data_out = 8'h9D;
                    16'hB3EB: data_out = 8'h9E;
                    16'hB3EC: data_out = 8'h9F;
                    16'hB3ED: data_out = 8'hA0;
                    16'hB3EE: data_out = 8'hA1;
                    16'hB3EF: data_out = 8'hA2;
                    16'hB3F0: data_out = 8'hA3;
                    16'hB3F1: data_out = 8'hA4;
                    16'hB3F2: data_out = 8'hA5;
                    16'hB3F3: data_out = 8'hA6;
                    16'hB3F4: data_out = 8'hA7;
                    16'hB3F5: data_out = 8'hA8;
                    16'hB3F6: data_out = 8'hA9;
                    16'hB3F7: data_out = 8'hAA;
                    16'hB3F8: data_out = 8'hAB;
                    16'hB3F9: data_out = 8'hAC;
                    16'hB3FA: data_out = 8'hAD;
                    16'hB3FB: data_out = 8'hAE;
                    16'hB3FC: data_out = 8'hAF;
                    16'hB3FD: data_out = 8'hB0;
                    16'hB3FE: data_out = 8'hB1;
                    16'hB3FF: data_out = 8'hB2;
                    16'hB400: data_out = 8'hB4;
                    16'hB401: data_out = 8'hB3;
                    16'hB402: data_out = 8'hB2;
                    16'hB403: data_out = 8'hB1;
                    16'hB404: data_out = 8'hB0;
                    16'hB405: data_out = 8'hAF;
                    16'hB406: data_out = 8'hAE;
                    16'hB407: data_out = 8'hAD;
                    16'hB408: data_out = 8'hAC;
                    16'hB409: data_out = 8'hAB;
                    16'hB40A: data_out = 8'hAA;
                    16'hB40B: data_out = 8'hA9;
                    16'hB40C: data_out = 8'hA8;
                    16'hB40D: data_out = 8'hA7;
                    16'hB40E: data_out = 8'hA6;
                    16'hB40F: data_out = 8'hA5;
                    16'hB410: data_out = 8'hA4;
                    16'hB411: data_out = 8'hA3;
                    16'hB412: data_out = 8'hA2;
                    16'hB413: data_out = 8'hA1;
                    16'hB414: data_out = 8'hA0;
                    16'hB415: data_out = 8'h9F;
                    16'hB416: data_out = 8'h9E;
                    16'hB417: data_out = 8'h9D;
                    16'hB418: data_out = 8'h9C;
                    16'hB419: data_out = 8'h9B;
                    16'hB41A: data_out = 8'h9A;
                    16'hB41B: data_out = 8'h99;
                    16'hB41C: data_out = 8'h98;
                    16'hB41D: data_out = 8'h97;
                    16'hB41E: data_out = 8'h96;
                    16'hB41F: data_out = 8'h95;
                    16'hB420: data_out = 8'h94;
                    16'hB421: data_out = 8'h93;
                    16'hB422: data_out = 8'h92;
                    16'hB423: data_out = 8'h91;
                    16'hB424: data_out = 8'h90;
                    16'hB425: data_out = 8'h8F;
                    16'hB426: data_out = 8'h8E;
                    16'hB427: data_out = 8'h8D;
                    16'hB428: data_out = 8'h8C;
                    16'hB429: data_out = 8'h8B;
                    16'hB42A: data_out = 8'h8A;
                    16'hB42B: data_out = 8'h89;
                    16'hB42C: data_out = 8'h88;
                    16'hB42D: data_out = 8'h87;
                    16'hB42E: data_out = 8'h86;
                    16'hB42F: data_out = 8'h85;
                    16'hB430: data_out = 8'h84;
                    16'hB431: data_out = 8'h83;
                    16'hB432: data_out = 8'h82;
                    16'hB433: data_out = 8'h81;
                    16'hB434: data_out = 8'h0;
                    16'hB435: data_out = 8'h1;
                    16'hB436: data_out = 8'h2;
                    16'hB437: data_out = 8'h3;
                    16'hB438: data_out = 8'h4;
                    16'hB439: data_out = 8'h5;
                    16'hB43A: data_out = 8'h6;
                    16'hB43B: data_out = 8'h7;
                    16'hB43C: data_out = 8'h8;
                    16'hB43D: data_out = 8'h9;
                    16'hB43E: data_out = 8'hA;
                    16'hB43F: data_out = 8'hB;
                    16'hB440: data_out = 8'hC;
                    16'hB441: data_out = 8'hD;
                    16'hB442: data_out = 8'hE;
                    16'hB443: data_out = 8'hF;
                    16'hB444: data_out = 8'h10;
                    16'hB445: data_out = 8'h11;
                    16'hB446: data_out = 8'h12;
                    16'hB447: data_out = 8'h13;
                    16'hB448: data_out = 8'h14;
                    16'hB449: data_out = 8'h15;
                    16'hB44A: data_out = 8'h16;
                    16'hB44B: data_out = 8'h17;
                    16'hB44C: data_out = 8'h18;
                    16'hB44D: data_out = 8'h19;
                    16'hB44E: data_out = 8'h1A;
                    16'hB44F: data_out = 8'h1B;
                    16'hB450: data_out = 8'h1C;
                    16'hB451: data_out = 8'h1D;
                    16'hB452: data_out = 8'h1E;
                    16'hB453: data_out = 8'h1F;
                    16'hB454: data_out = 8'h20;
                    16'hB455: data_out = 8'h21;
                    16'hB456: data_out = 8'h22;
                    16'hB457: data_out = 8'h23;
                    16'hB458: data_out = 8'h24;
                    16'hB459: data_out = 8'h25;
                    16'hB45A: data_out = 8'h26;
                    16'hB45B: data_out = 8'h27;
                    16'hB45C: data_out = 8'h28;
                    16'hB45D: data_out = 8'h29;
                    16'hB45E: data_out = 8'h2A;
                    16'hB45F: data_out = 8'h2B;
                    16'hB460: data_out = 8'h2C;
                    16'hB461: data_out = 8'h2D;
                    16'hB462: data_out = 8'h2E;
                    16'hB463: data_out = 8'h2F;
                    16'hB464: data_out = 8'h30;
                    16'hB465: data_out = 8'h31;
                    16'hB466: data_out = 8'h32;
                    16'hB467: data_out = 8'h33;
                    16'hB468: data_out = 8'h34;
                    16'hB469: data_out = 8'h35;
                    16'hB46A: data_out = 8'h36;
                    16'hB46B: data_out = 8'h37;
                    16'hB46C: data_out = 8'h38;
                    16'hB46D: data_out = 8'h39;
                    16'hB46E: data_out = 8'h3A;
                    16'hB46F: data_out = 8'h3B;
                    16'hB470: data_out = 8'h3C;
                    16'hB471: data_out = 8'h3D;
                    16'hB472: data_out = 8'h3E;
                    16'hB473: data_out = 8'h3F;
                    16'hB474: data_out = 8'h40;
                    16'hB475: data_out = 8'h41;
                    16'hB476: data_out = 8'h42;
                    16'hB477: data_out = 8'h43;
                    16'hB478: data_out = 8'h44;
                    16'hB479: data_out = 8'h45;
                    16'hB47A: data_out = 8'h46;
                    16'hB47B: data_out = 8'h47;
                    16'hB47C: data_out = 8'h48;
                    16'hB47D: data_out = 8'h49;
                    16'hB47E: data_out = 8'h4A;
                    16'hB47F: data_out = 8'h4B;
                    16'hB480: data_out = 8'hB4;
                    16'hB481: data_out = 8'hB5;
                    16'hB482: data_out = 8'hB6;
                    16'hB483: data_out = 8'hB7;
                    16'hB484: data_out = 8'hB8;
                    16'hB485: data_out = 8'hB9;
                    16'hB486: data_out = 8'hBA;
                    16'hB487: data_out = 8'hBB;
                    16'hB488: data_out = 8'hBC;
                    16'hB489: data_out = 8'hBD;
                    16'hB48A: data_out = 8'hBE;
                    16'hB48B: data_out = 8'hBF;
                    16'hB48C: data_out = 8'hC0;
                    16'hB48D: data_out = 8'hC1;
                    16'hB48E: data_out = 8'hC2;
                    16'hB48F: data_out = 8'hC3;
                    16'hB490: data_out = 8'hC4;
                    16'hB491: data_out = 8'hC5;
                    16'hB492: data_out = 8'hC6;
                    16'hB493: data_out = 8'hC7;
                    16'hB494: data_out = 8'hC8;
                    16'hB495: data_out = 8'hC9;
                    16'hB496: data_out = 8'hCA;
                    16'hB497: data_out = 8'hCB;
                    16'hB498: data_out = 8'hCC;
                    16'hB499: data_out = 8'hCD;
                    16'hB49A: data_out = 8'hCE;
                    16'hB49B: data_out = 8'hCF;
                    16'hB49C: data_out = 8'hD0;
                    16'hB49D: data_out = 8'hD1;
                    16'hB49E: data_out = 8'hD2;
                    16'hB49F: data_out = 8'hD3;
                    16'hB4A0: data_out = 8'hD4;
                    16'hB4A1: data_out = 8'hD5;
                    16'hB4A2: data_out = 8'hD6;
                    16'hB4A3: data_out = 8'hD7;
                    16'hB4A4: data_out = 8'hD8;
                    16'hB4A5: data_out = 8'hD9;
                    16'hB4A6: data_out = 8'hDA;
                    16'hB4A7: data_out = 8'hDB;
                    16'hB4A8: data_out = 8'hDC;
                    16'hB4A9: data_out = 8'hDD;
                    16'hB4AA: data_out = 8'hDE;
                    16'hB4AB: data_out = 8'hDF;
                    16'hB4AC: data_out = 8'hE0;
                    16'hB4AD: data_out = 8'hE1;
                    16'hB4AE: data_out = 8'hE2;
                    16'hB4AF: data_out = 8'hE3;
                    16'hB4B0: data_out = 8'hE4;
                    16'hB4B1: data_out = 8'hE5;
                    16'hB4B2: data_out = 8'hE6;
                    16'hB4B3: data_out = 8'hE7;
                    16'hB4B4: data_out = 8'hE8;
                    16'hB4B5: data_out = 8'hE9;
                    16'hB4B6: data_out = 8'hEA;
                    16'hB4B7: data_out = 8'hEB;
                    16'hB4B8: data_out = 8'hEC;
                    16'hB4B9: data_out = 8'hED;
                    16'hB4BA: data_out = 8'hEE;
                    16'hB4BB: data_out = 8'hEF;
                    16'hB4BC: data_out = 8'hF0;
                    16'hB4BD: data_out = 8'hF1;
                    16'hB4BE: data_out = 8'hF2;
                    16'hB4BF: data_out = 8'hF3;
                    16'hB4C0: data_out = 8'hF4;
                    16'hB4C1: data_out = 8'hF5;
                    16'hB4C2: data_out = 8'hF6;
                    16'hB4C3: data_out = 8'hF7;
                    16'hB4C4: data_out = 8'hF8;
                    16'hB4C5: data_out = 8'hF9;
                    16'hB4C6: data_out = 8'hFA;
                    16'hB4C7: data_out = 8'hFB;
                    16'hB4C8: data_out = 8'hFC;
                    16'hB4C9: data_out = 8'hFD;
                    16'hB4CA: data_out = 8'hFE;
                    16'hB4CB: data_out = 8'hFF;
                    16'hB4CC: data_out = 8'h80;
                    16'hB4CD: data_out = 8'h81;
                    16'hB4CE: data_out = 8'h82;
                    16'hB4CF: data_out = 8'h83;
                    16'hB4D0: data_out = 8'h84;
                    16'hB4D1: data_out = 8'h85;
                    16'hB4D2: data_out = 8'h86;
                    16'hB4D3: data_out = 8'h87;
                    16'hB4D4: data_out = 8'h88;
                    16'hB4D5: data_out = 8'h89;
                    16'hB4D6: data_out = 8'h8A;
                    16'hB4D7: data_out = 8'h8B;
                    16'hB4D8: data_out = 8'h8C;
                    16'hB4D9: data_out = 8'h8D;
                    16'hB4DA: data_out = 8'h8E;
                    16'hB4DB: data_out = 8'h8F;
                    16'hB4DC: data_out = 8'h90;
                    16'hB4DD: data_out = 8'h91;
                    16'hB4DE: data_out = 8'h92;
                    16'hB4DF: data_out = 8'h93;
                    16'hB4E0: data_out = 8'h94;
                    16'hB4E1: data_out = 8'h95;
                    16'hB4E2: data_out = 8'h96;
                    16'hB4E3: data_out = 8'h97;
                    16'hB4E4: data_out = 8'h98;
                    16'hB4E5: data_out = 8'h99;
                    16'hB4E6: data_out = 8'h9A;
                    16'hB4E7: data_out = 8'h9B;
                    16'hB4E8: data_out = 8'h9C;
                    16'hB4E9: data_out = 8'h9D;
                    16'hB4EA: data_out = 8'h9E;
                    16'hB4EB: data_out = 8'h9F;
                    16'hB4EC: data_out = 8'hA0;
                    16'hB4ED: data_out = 8'hA1;
                    16'hB4EE: data_out = 8'hA2;
                    16'hB4EF: data_out = 8'hA3;
                    16'hB4F0: data_out = 8'hA4;
                    16'hB4F1: data_out = 8'hA5;
                    16'hB4F2: data_out = 8'hA6;
                    16'hB4F3: data_out = 8'hA7;
                    16'hB4F4: data_out = 8'hA8;
                    16'hB4F5: data_out = 8'hA9;
                    16'hB4F6: data_out = 8'hAA;
                    16'hB4F7: data_out = 8'hAB;
                    16'hB4F8: data_out = 8'hAC;
                    16'hB4F9: data_out = 8'hAD;
                    16'hB4FA: data_out = 8'hAE;
                    16'hB4FB: data_out = 8'hAF;
                    16'hB4FC: data_out = 8'hB0;
                    16'hB4FD: data_out = 8'hB1;
                    16'hB4FE: data_out = 8'hB2;
                    16'hB4FF: data_out = 8'hB3;
                    16'hB500: data_out = 8'hB5;
                    16'hB501: data_out = 8'hB4;
                    16'hB502: data_out = 8'hB3;
                    16'hB503: data_out = 8'hB2;
                    16'hB504: data_out = 8'hB1;
                    16'hB505: data_out = 8'hB0;
                    16'hB506: data_out = 8'hAF;
                    16'hB507: data_out = 8'hAE;
                    16'hB508: data_out = 8'hAD;
                    16'hB509: data_out = 8'hAC;
                    16'hB50A: data_out = 8'hAB;
                    16'hB50B: data_out = 8'hAA;
                    16'hB50C: data_out = 8'hA9;
                    16'hB50D: data_out = 8'hA8;
                    16'hB50E: data_out = 8'hA7;
                    16'hB50F: data_out = 8'hA6;
                    16'hB510: data_out = 8'hA5;
                    16'hB511: data_out = 8'hA4;
                    16'hB512: data_out = 8'hA3;
                    16'hB513: data_out = 8'hA2;
                    16'hB514: data_out = 8'hA1;
                    16'hB515: data_out = 8'hA0;
                    16'hB516: data_out = 8'h9F;
                    16'hB517: data_out = 8'h9E;
                    16'hB518: data_out = 8'h9D;
                    16'hB519: data_out = 8'h9C;
                    16'hB51A: data_out = 8'h9B;
                    16'hB51B: data_out = 8'h9A;
                    16'hB51C: data_out = 8'h99;
                    16'hB51D: data_out = 8'h98;
                    16'hB51E: data_out = 8'h97;
                    16'hB51F: data_out = 8'h96;
                    16'hB520: data_out = 8'h95;
                    16'hB521: data_out = 8'h94;
                    16'hB522: data_out = 8'h93;
                    16'hB523: data_out = 8'h92;
                    16'hB524: data_out = 8'h91;
                    16'hB525: data_out = 8'h90;
                    16'hB526: data_out = 8'h8F;
                    16'hB527: data_out = 8'h8E;
                    16'hB528: data_out = 8'h8D;
                    16'hB529: data_out = 8'h8C;
                    16'hB52A: data_out = 8'h8B;
                    16'hB52B: data_out = 8'h8A;
                    16'hB52C: data_out = 8'h89;
                    16'hB52D: data_out = 8'h88;
                    16'hB52E: data_out = 8'h87;
                    16'hB52F: data_out = 8'h86;
                    16'hB530: data_out = 8'h85;
                    16'hB531: data_out = 8'h84;
                    16'hB532: data_out = 8'h83;
                    16'hB533: data_out = 8'h82;
                    16'hB534: data_out = 8'h81;
                    16'hB535: data_out = 8'h0;
                    16'hB536: data_out = 8'h1;
                    16'hB537: data_out = 8'h2;
                    16'hB538: data_out = 8'h3;
                    16'hB539: data_out = 8'h4;
                    16'hB53A: data_out = 8'h5;
                    16'hB53B: data_out = 8'h6;
                    16'hB53C: data_out = 8'h7;
                    16'hB53D: data_out = 8'h8;
                    16'hB53E: data_out = 8'h9;
                    16'hB53F: data_out = 8'hA;
                    16'hB540: data_out = 8'hB;
                    16'hB541: data_out = 8'hC;
                    16'hB542: data_out = 8'hD;
                    16'hB543: data_out = 8'hE;
                    16'hB544: data_out = 8'hF;
                    16'hB545: data_out = 8'h10;
                    16'hB546: data_out = 8'h11;
                    16'hB547: data_out = 8'h12;
                    16'hB548: data_out = 8'h13;
                    16'hB549: data_out = 8'h14;
                    16'hB54A: data_out = 8'h15;
                    16'hB54B: data_out = 8'h16;
                    16'hB54C: data_out = 8'h17;
                    16'hB54D: data_out = 8'h18;
                    16'hB54E: data_out = 8'h19;
                    16'hB54F: data_out = 8'h1A;
                    16'hB550: data_out = 8'h1B;
                    16'hB551: data_out = 8'h1C;
                    16'hB552: data_out = 8'h1D;
                    16'hB553: data_out = 8'h1E;
                    16'hB554: data_out = 8'h1F;
                    16'hB555: data_out = 8'h20;
                    16'hB556: data_out = 8'h21;
                    16'hB557: data_out = 8'h22;
                    16'hB558: data_out = 8'h23;
                    16'hB559: data_out = 8'h24;
                    16'hB55A: data_out = 8'h25;
                    16'hB55B: data_out = 8'h26;
                    16'hB55C: data_out = 8'h27;
                    16'hB55D: data_out = 8'h28;
                    16'hB55E: data_out = 8'h29;
                    16'hB55F: data_out = 8'h2A;
                    16'hB560: data_out = 8'h2B;
                    16'hB561: data_out = 8'h2C;
                    16'hB562: data_out = 8'h2D;
                    16'hB563: data_out = 8'h2E;
                    16'hB564: data_out = 8'h2F;
                    16'hB565: data_out = 8'h30;
                    16'hB566: data_out = 8'h31;
                    16'hB567: data_out = 8'h32;
                    16'hB568: data_out = 8'h33;
                    16'hB569: data_out = 8'h34;
                    16'hB56A: data_out = 8'h35;
                    16'hB56B: data_out = 8'h36;
                    16'hB56C: data_out = 8'h37;
                    16'hB56D: data_out = 8'h38;
                    16'hB56E: data_out = 8'h39;
                    16'hB56F: data_out = 8'h3A;
                    16'hB570: data_out = 8'h3B;
                    16'hB571: data_out = 8'h3C;
                    16'hB572: data_out = 8'h3D;
                    16'hB573: data_out = 8'h3E;
                    16'hB574: data_out = 8'h3F;
                    16'hB575: data_out = 8'h40;
                    16'hB576: data_out = 8'h41;
                    16'hB577: data_out = 8'h42;
                    16'hB578: data_out = 8'h43;
                    16'hB579: data_out = 8'h44;
                    16'hB57A: data_out = 8'h45;
                    16'hB57B: data_out = 8'h46;
                    16'hB57C: data_out = 8'h47;
                    16'hB57D: data_out = 8'h48;
                    16'hB57E: data_out = 8'h49;
                    16'hB57F: data_out = 8'h4A;
                    16'hB580: data_out = 8'hB5;
                    16'hB581: data_out = 8'hB6;
                    16'hB582: data_out = 8'hB7;
                    16'hB583: data_out = 8'hB8;
                    16'hB584: data_out = 8'hB9;
                    16'hB585: data_out = 8'hBA;
                    16'hB586: data_out = 8'hBB;
                    16'hB587: data_out = 8'hBC;
                    16'hB588: data_out = 8'hBD;
                    16'hB589: data_out = 8'hBE;
                    16'hB58A: data_out = 8'hBF;
                    16'hB58B: data_out = 8'hC0;
                    16'hB58C: data_out = 8'hC1;
                    16'hB58D: data_out = 8'hC2;
                    16'hB58E: data_out = 8'hC3;
                    16'hB58F: data_out = 8'hC4;
                    16'hB590: data_out = 8'hC5;
                    16'hB591: data_out = 8'hC6;
                    16'hB592: data_out = 8'hC7;
                    16'hB593: data_out = 8'hC8;
                    16'hB594: data_out = 8'hC9;
                    16'hB595: data_out = 8'hCA;
                    16'hB596: data_out = 8'hCB;
                    16'hB597: data_out = 8'hCC;
                    16'hB598: data_out = 8'hCD;
                    16'hB599: data_out = 8'hCE;
                    16'hB59A: data_out = 8'hCF;
                    16'hB59B: data_out = 8'hD0;
                    16'hB59C: data_out = 8'hD1;
                    16'hB59D: data_out = 8'hD2;
                    16'hB59E: data_out = 8'hD3;
                    16'hB59F: data_out = 8'hD4;
                    16'hB5A0: data_out = 8'hD5;
                    16'hB5A1: data_out = 8'hD6;
                    16'hB5A2: data_out = 8'hD7;
                    16'hB5A3: data_out = 8'hD8;
                    16'hB5A4: data_out = 8'hD9;
                    16'hB5A5: data_out = 8'hDA;
                    16'hB5A6: data_out = 8'hDB;
                    16'hB5A7: data_out = 8'hDC;
                    16'hB5A8: data_out = 8'hDD;
                    16'hB5A9: data_out = 8'hDE;
                    16'hB5AA: data_out = 8'hDF;
                    16'hB5AB: data_out = 8'hE0;
                    16'hB5AC: data_out = 8'hE1;
                    16'hB5AD: data_out = 8'hE2;
                    16'hB5AE: data_out = 8'hE3;
                    16'hB5AF: data_out = 8'hE4;
                    16'hB5B0: data_out = 8'hE5;
                    16'hB5B1: data_out = 8'hE6;
                    16'hB5B2: data_out = 8'hE7;
                    16'hB5B3: data_out = 8'hE8;
                    16'hB5B4: data_out = 8'hE9;
                    16'hB5B5: data_out = 8'hEA;
                    16'hB5B6: data_out = 8'hEB;
                    16'hB5B7: data_out = 8'hEC;
                    16'hB5B8: data_out = 8'hED;
                    16'hB5B9: data_out = 8'hEE;
                    16'hB5BA: data_out = 8'hEF;
                    16'hB5BB: data_out = 8'hF0;
                    16'hB5BC: data_out = 8'hF1;
                    16'hB5BD: data_out = 8'hF2;
                    16'hB5BE: data_out = 8'hF3;
                    16'hB5BF: data_out = 8'hF4;
                    16'hB5C0: data_out = 8'hF5;
                    16'hB5C1: data_out = 8'hF6;
                    16'hB5C2: data_out = 8'hF7;
                    16'hB5C3: data_out = 8'hF8;
                    16'hB5C4: data_out = 8'hF9;
                    16'hB5C5: data_out = 8'hFA;
                    16'hB5C6: data_out = 8'hFB;
                    16'hB5C7: data_out = 8'hFC;
                    16'hB5C8: data_out = 8'hFD;
                    16'hB5C9: data_out = 8'hFE;
                    16'hB5CA: data_out = 8'hFF;
                    16'hB5CB: data_out = 8'h80;
                    16'hB5CC: data_out = 8'h81;
                    16'hB5CD: data_out = 8'h82;
                    16'hB5CE: data_out = 8'h83;
                    16'hB5CF: data_out = 8'h84;
                    16'hB5D0: data_out = 8'h85;
                    16'hB5D1: data_out = 8'h86;
                    16'hB5D2: data_out = 8'h87;
                    16'hB5D3: data_out = 8'h88;
                    16'hB5D4: data_out = 8'h89;
                    16'hB5D5: data_out = 8'h8A;
                    16'hB5D6: data_out = 8'h8B;
                    16'hB5D7: data_out = 8'h8C;
                    16'hB5D8: data_out = 8'h8D;
                    16'hB5D9: data_out = 8'h8E;
                    16'hB5DA: data_out = 8'h8F;
                    16'hB5DB: data_out = 8'h90;
                    16'hB5DC: data_out = 8'h91;
                    16'hB5DD: data_out = 8'h92;
                    16'hB5DE: data_out = 8'h93;
                    16'hB5DF: data_out = 8'h94;
                    16'hB5E0: data_out = 8'h95;
                    16'hB5E1: data_out = 8'h96;
                    16'hB5E2: data_out = 8'h97;
                    16'hB5E3: data_out = 8'h98;
                    16'hB5E4: data_out = 8'h99;
                    16'hB5E5: data_out = 8'h9A;
                    16'hB5E6: data_out = 8'h9B;
                    16'hB5E7: data_out = 8'h9C;
                    16'hB5E8: data_out = 8'h9D;
                    16'hB5E9: data_out = 8'h9E;
                    16'hB5EA: data_out = 8'h9F;
                    16'hB5EB: data_out = 8'hA0;
                    16'hB5EC: data_out = 8'hA1;
                    16'hB5ED: data_out = 8'hA2;
                    16'hB5EE: data_out = 8'hA3;
                    16'hB5EF: data_out = 8'hA4;
                    16'hB5F0: data_out = 8'hA5;
                    16'hB5F1: data_out = 8'hA6;
                    16'hB5F2: data_out = 8'hA7;
                    16'hB5F3: data_out = 8'hA8;
                    16'hB5F4: data_out = 8'hA9;
                    16'hB5F5: data_out = 8'hAA;
                    16'hB5F6: data_out = 8'hAB;
                    16'hB5F7: data_out = 8'hAC;
                    16'hB5F8: data_out = 8'hAD;
                    16'hB5F9: data_out = 8'hAE;
                    16'hB5FA: data_out = 8'hAF;
                    16'hB5FB: data_out = 8'hB0;
                    16'hB5FC: data_out = 8'hB1;
                    16'hB5FD: data_out = 8'hB2;
                    16'hB5FE: data_out = 8'hB3;
                    16'hB5FF: data_out = 8'hB4;
                    16'hB600: data_out = 8'hB6;
                    16'hB601: data_out = 8'hB5;
                    16'hB602: data_out = 8'hB4;
                    16'hB603: data_out = 8'hB3;
                    16'hB604: data_out = 8'hB2;
                    16'hB605: data_out = 8'hB1;
                    16'hB606: data_out = 8'hB0;
                    16'hB607: data_out = 8'hAF;
                    16'hB608: data_out = 8'hAE;
                    16'hB609: data_out = 8'hAD;
                    16'hB60A: data_out = 8'hAC;
                    16'hB60B: data_out = 8'hAB;
                    16'hB60C: data_out = 8'hAA;
                    16'hB60D: data_out = 8'hA9;
                    16'hB60E: data_out = 8'hA8;
                    16'hB60F: data_out = 8'hA7;
                    16'hB610: data_out = 8'hA6;
                    16'hB611: data_out = 8'hA5;
                    16'hB612: data_out = 8'hA4;
                    16'hB613: data_out = 8'hA3;
                    16'hB614: data_out = 8'hA2;
                    16'hB615: data_out = 8'hA1;
                    16'hB616: data_out = 8'hA0;
                    16'hB617: data_out = 8'h9F;
                    16'hB618: data_out = 8'h9E;
                    16'hB619: data_out = 8'h9D;
                    16'hB61A: data_out = 8'h9C;
                    16'hB61B: data_out = 8'h9B;
                    16'hB61C: data_out = 8'h9A;
                    16'hB61D: data_out = 8'h99;
                    16'hB61E: data_out = 8'h98;
                    16'hB61F: data_out = 8'h97;
                    16'hB620: data_out = 8'h96;
                    16'hB621: data_out = 8'h95;
                    16'hB622: data_out = 8'h94;
                    16'hB623: data_out = 8'h93;
                    16'hB624: data_out = 8'h92;
                    16'hB625: data_out = 8'h91;
                    16'hB626: data_out = 8'h90;
                    16'hB627: data_out = 8'h8F;
                    16'hB628: data_out = 8'h8E;
                    16'hB629: data_out = 8'h8D;
                    16'hB62A: data_out = 8'h8C;
                    16'hB62B: data_out = 8'h8B;
                    16'hB62C: data_out = 8'h8A;
                    16'hB62D: data_out = 8'h89;
                    16'hB62E: data_out = 8'h88;
                    16'hB62F: data_out = 8'h87;
                    16'hB630: data_out = 8'h86;
                    16'hB631: data_out = 8'h85;
                    16'hB632: data_out = 8'h84;
                    16'hB633: data_out = 8'h83;
                    16'hB634: data_out = 8'h82;
                    16'hB635: data_out = 8'h81;
                    16'hB636: data_out = 8'h0;
                    16'hB637: data_out = 8'h1;
                    16'hB638: data_out = 8'h2;
                    16'hB639: data_out = 8'h3;
                    16'hB63A: data_out = 8'h4;
                    16'hB63B: data_out = 8'h5;
                    16'hB63C: data_out = 8'h6;
                    16'hB63D: data_out = 8'h7;
                    16'hB63E: data_out = 8'h8;
                    16'hB63F: data_out = 8'h9;
                    16'hB640: data_out = 8'hA;
                    16'hB641: data_out = 8'hB;
                    16'hB642: data_out = 8'hC;
                    16'hB643: data_out = 8'hD;
                    16'hB644: data_out = 8'hE;
                    16'hB645: data_out = 8'hF;
                    16'hB646: data_out = 8'h10;
                    16'hB647: data_out = 8'h11;
                    16'hB648: data_out = 8'h12;
                    16'hB649: data_out = 8'h13;
                    16'hB64A: data_out = 8'h14;
                    16'hB64B: data_out = 8'h15;
                    16'hB64C: data_out = 8'h16;
                    16'hB64D: data_out = 8'h17;
                    16'hB64E: data_out = 8'h18;
                    16'hB64F: data_out = 8'h19;
                    16'hB650: data_out = 8'h1A;
                    16'hB651: data_out = 8'h1B;
                    16'hB652: data_out = 8'h1C;
                    16'hB653: data_out = 8'h1D;
                    16'hB654: data_out = 8'h1E;
                    16'hB655: data_out = 8'h1F;
                    16'hB656: data_out = 8'h20;
                    16'hB657: data_out = 8'h21;
                    16'hB658: data_out = 8'h22;
                    16'hB659: data_out = 8'h23;
                    16'hB65A: data_out = 8'h24;
                    16'hB65B: data_out = 8'h25;
                    16'hB65C: data_out = 8'h26;
                    16'hB65D: data_out = 8'h27;
                    16'hB65E: data_out = 8'h28;
                    16'hB65F: data_out = 8'h29;
                    16'hB660: data_out = 8'h2A;
                    16'hB661: data_out = 8'h2B;
                    16'hB662: data_out = 8'h2C;
                    16'hB663: data_out = 8'h2D;
                    16'hB664: data_out = 8'h2E;
                    16'hB665: data_out = 8'h2F;
                    16'hB666: data_out = 8'h30;
                    16'hB667: data_out = 8'h31;
                    16'hB668: data_out = 8'h32;
                    16'hB669: data_out = 8'h33;
                    16'hB66A: data_out = 8'h34;
                    16'hB66B: data_out = 8'h35;
                    16'hB66C: data_out = 8'h36;
                    16'hB66D: data_out = 8'h37;
                    16'hB66E: data_out = 8'h38;
                    16'hB66F: data_out = 8'h39;
                    16'hB670: data_out = 8'h3A;
                    16'hB671: data_out = 8'h3B;
                    16'hB672: data_out = 8'h3C;
                    16'hB673: data_out = 8'h3D;
                    16'hB674: data_out = 8'h3E;
                    16'hB675: data_out = 8'h3F;
                    16'hB676: data_out = 8'h40;
                    16'hB677: data_out = 8'h41;
                    16'hB678: data_out = 8'h42;
                    16'hB679: data_out = 8'h43;
                    16'hB67A: data_out = 8'h44;
                    16'hB67B: data_out = 8'h45;
                    16'hB67C: data_out = 8'h46;
                    16'hB67D: data_out = 8'h47;
                    16'hB67E: data_out = 8'h48;
                    16'hB67F: data_out = 8'h49;
                    16'hB680: data_out = 8'hB6;
                    16'hB681: data_out = 8'hB7;
                    16'hB682: data_out = 8'hB8;
                    16'hB683: data_out = 8'hB9;
                    16'hB684: data_out = 8'hBA;
                    16'hB685: data_out = 8'hBB;
                    16'hB686: data_out = 8'hBC;
                    16'hB687: data_out = 8'hBD;
                    16'hB688: data_out = 8'hBE;
                    16'hB689: data_out = 8'hBF;
                    16'hB68A: data_out = 8'hC0;
                    16'hB68B: data_out = 8'hC1;
                    16'hB68C: data_out = 8'hC2;
                    16'hB68D: data_out = 8'hC3;
                    16'hB68E: data_out = 8'hC4;
                    16'hB68F: data_out = 8'hC5;
                    16'hB690: data_out = 8'hC6;
                    16'hB691: data_out = 8'hC7;
                    16'hB692: data_out = 8'hC8;
                    16'hB693: data_out = 8'hC9;
                    16'hB694: data_out = 8'hCA;
                    16'hB695: data_out = 8'hCB;
                    16'hB696: data_out = 8'hCC;
                    16'hB697: data_out = 8'hCD;
                    16'hB698: data_out = 8'hCE;
                    16'hB699: data_out = 8'hCF;
                    16'hB69A: data_out = 8'hD0;
                    16'hB69B: data_out = 8'hD1;
                    16'hB69C: data_out = 8'hD2;
                    16'hB69D: data_out = 8'hD3;
                    16'hB69E: data_out = 8'hD4;
                    16'hB69F: data_out = 8'hD5;
                    16'hB6A0: data_out = 8'hD6;
                    16'hB6A1: data_out = 8'hD7;
                    16'hB6A2: data_out = 8'hD8;
                    16'hB6A3: data_out = 8'hD9;
                    16'hB6A4: data_out = 8'hDA;
                    16'hB6A5: data_out = 8'hDB;
                    16'hB6A6: data_out = 8'hDC;
                    16'hB6A7: data_out = 8'hDD;
                    16'hB6A8: data_out = 8'hDE;
                    16'hB6A9: data_out = 8'hDF;
                    16'hB6AA: data_out = 8'hE0;
                    16'hB6AB: data_out = 8'hE1;
                    16'hB6AC: data_out = 8'hE2;
                    16'hB6AD: data_out = 8'hE3;
                    16'hB6AE: data_out = 8'hE4;
                    16'hB6AF: data_out = 8'hE5;
                    16'hB6B0: data_out = 8'hE6;
                    16'hB6B1: data_out = 8'hE7;
                    16'hB6B2: data_out = 8'hE8;
                    16'hB6B3: data_out = 8'hE9;
                    16'hB6B4: data_out = 8'hEA;
                    16'hB6B5: data_out = 8'hEB;
                    16'hB6B6: data_out = 8'hEC;
                    16'hB6B7: data_out = 8'hED;
                    16'hB6B8: data_out = 8'hEE;
                    16'hB6B9: data_out = 8'hEF;
                    16'hB6BA: data_out = 8'hF0;
                    16'hB6BB: data_out = 8'hF1;
                    16'hB6BC: data_out = 8'hF2;
                    16'hB6BD: data_out = 8'hF3;
                    16'hB6BE: data_out = 8'hF4;
                    16'hB6BF: data_out = 8'hF5;
                    16'hB6C0: data_out = 8'hF6;
                    16'hB6C1: data_out = 8'hF7;
                    16'hB6C2: data_out = 8'hF8;
                    16'hB6C3: data_out = 8'hF9;
                    16'hB6C4: data_out = 8'hFA;
                    16'hB6C5: data_out = 8'hFB;
                    16'hB6C6: data_out = 8'hFC;
                    16'hB6C7: data_out = 8'hFD;
                    16'hB6C8: data_out = 8'hFE;
                    16'hB6C9: data_out = 8'hFF;
                    16'hB6CA: data_out = 8'h80;
                    16'hB6CB: data_out = 8'h81;
                    16'hB6CC: data_out = 8'h82;
                    16'hB6CD: data_out = 8'h83;
                    16'hB6CE: data_out = 8'h84;
                    16'hB6CF: data_out = 8'h85;
                    16'hB6D0: data_out = 8'h86;
                    16'hB6D1: data_out = 8'h87;
                    16'hB6D2: data_out = 8'h88;
                    16'hB6D3: data_out = 8'h89;
                    16'hB6D4: data_out = 8'h8A;
                    16'hB6D5: data_out = 8'h8B;
                    16'hB6D6: data_out = 8'h8C;
                    16'hB6D7: data_out = 8'h8D;
                    16'hB6D8: data_out = 8'h8E;
                    16'hB6D9: data_out = 8'h8F;
                    16'hB6DA: data_out = 8'h90;
                    16'hB6DB: data_out = 8'h91;
                    16'hB6DC: data_out = 8'h92;
                    16'hB6DD: data_out = 8'h93;
                    16'hB6DE: data_out = 8'h94;
                    16'hB6DF: data_out = 8'h95;
                    16'hB6E0: data_out = 8'h96;
                    16'hB6E1: data_out = 8'h97;
                    16'hB6E2: data_out = 8'h98;
                    16'hB6E3: data_out = 8'h99;
                    16'hB6E4: data_out = 8'h9A;
                    16'hB6E5: data_out = 8'h9B;
                    16'hB6E6: data_out = 8'h9C;
                    16'hB6E7: data_out = 8'h9D;
                    16'hB6E8: data_out = 8'h9E;
                    16'hB6E9: data_out = 8'h9F;
                    16'hB6EA: data_out = 8'hA0;
                    16'hB6EB: data_out = 8'hA1;
                    16'hB6EC: data_out = 8'hA2;
                    16'hB6ED: data_out = 8'hA3;
                    16'hB6EE: data_out = 8'hA4;
                    16'hB6EF: data_out = 8'hA5;
                    16'hB6F0: data_out = 8'hA6;
                    16'hB6F1: data_out = 8'hA7;
                    16'hB6F2: data_out = 8'hA8;
                    16'hB6F3: data_out = 8'hA9;
                    16'hB6F4: data_out = 8'hAA;
                    16'hB6F5: data_out = 8'hAB;
                    16'hB6F6: data_out = 8'hAC;
                    16'hB6F7: data_out = 8'hAD;
                    16'hB6F8: data_out = 8'hAE;
                    16'hB6F9: data_out = 8'hAF;
                    16'hB6FA: data_out = 8'hB0;
                    16'hB6FB: data_out = 8'hB1;
                    16'hB6FC: data_out = 8'hB2;
                    16'hB6FD: data_out = 8'hB3;
                    16'hB6FE: data_out = 8'hB4;
                    16'hB6FF: data_out = 8'hB5;
                    16'hB700: data_out = 8'hB7;
                    16'hB701: data_out = 8'hB6;
                    16'hB702: data_out = 8'hB5;
                    16'hB703: data_out = 8'hB4;
                    16'hB704: data_out = 8'hB3;
                    16'hB705: data_out = 8'hB2;
                    16'hB706: data_out = 8'hB1;
                    16'hB707: data_out = 8'hB0;
                    16'hB708: data_out = 8'hAF;
                    16'hB709: data_out = 8'hAE;
                    16'hB70A: data_out = 8'hAD;
                    16'hB70B: data_out = 8'hAC;
                    16'hB70C: data_out = 8'hAB;
                    16'hB70D: data_out = 8'hAA;
                    16'hB70E: data_out = 8'hA9;
                    16'hB70F: data_out = 8'hA8;
                    16'hB710: data_out = 8'hA7;
                    16'hB711: data_out = 8'hA6;
                    16'hB712: data_out = 8'hA5;
                    16'hB713: data_out = 8'hA4;
                    16'hB714: data_out = 8'hA3;
                    16'hB715: data_out = 8'hA2;
                    16'hB716: data_out = 8'hA1;
                    16'hB717: data_out = 8'hA0;
                    16'hB718: data_out = 8'h9F;
                    16'hB719: data_out = 8'h9E;
                    16'hB71A: data_out = 8'h9D;
                    16'hB71B: data_out = 8'h9C;
                    16'hB71C: data_out = 8'h9B;
                    16'hB71D: data_out = 8'h9A;
                    16'hB71E: data_out = 8'h99;
                    16'hB71F: data_out = 8'h98;
                    16'hB720: data_out = 8'h97;
                    16'hB721: data_out = 8'h96;
                    16'hB722: data_out = 8'h95;
                    16'hB723: data_out = 8'h94;
                    16'hB724: data_out = 8'h93;
                    16'hB725: data_out = 8'h92;
                    16'hB726: data_out = 8'h91;
                    16'hB727: data_out = 8'h90;
                    16'hB728: data_out = 8'h8F;
                    16'hB729: data_out = 8'h8E;
                    16'hB72A: data_out = 8'h8D;
                    16'hB72B: data_out = 8'h8C;
                    16'hB72C: data_out = 8'h8B;
                    16'hB72D: data_out = 8'h8A;
                    16'hB72E: data_out = 8'h89;
                    16'hB72F: data_out = 8'h88;
                    16'hB730: data_out = 8'h87;
                    16'hB731: data_out = 8'h86;
                    16'hB732: data_out = 8'h85;
                    16'hB733: data_out = 8'h84;
                    16'hB734: data_out = 8'h83;
                    16'hB735: data_out = 8'h82;
                    16'hB736: data_out = 8'h81;
                    16'hB737: data_out = 8'h0;
                    16'hB738: data_out = 8'h1;
                    16'hB739: data_out = 8'h2;
                    16'hB73A: data_out = 8'h3;
                    16'hB73B: data_out = 8'h4;
                    16'hB73C: data_out = 8'h5;
                    16'hB73D: data_out = 8'h6;
                    16'hB73E: data_out = 8'h7;
                    16'hB73F: data_out = 8'h8;
                    16'hB740: data_out = 8'h9;
                    16'hB741: data_out = 8'hA;
                    16'hB742: data_out = 8'hB;
                    16'hB743: data_out = 8'hC;
                    16'hB744: data_out = 8'hD;
                    16'hB745: data_out = 8'hE;
                    16'hB746: data_out = 8'hF;
                    16'hB747: data_out = 8'h10;
                    16'hB748: data_out = 8'h11;
                    16'hB749: data_out = 8'h12;
                    16'hB74A: data_out = 8'h13;
                    16'hB74B: data_out = 8'h14;
                    16'hB74C: data_out = 8'h15;
                    16'hB74D: data_out = 8'h16;
                    16'hB74E: data_out = 8'h17;
                    16'hB74F: data_out = 8'h18;
                    16'hB750: data_out = 8'h19;
                    16'hB751: data_out = 8'h1A;
                    16'hB752: data_out = 8'h1B;
                    16'hB753: data_out = 8'h1C;
                    16'hB754: data_out = 8'h1D;
                    16'hB755: data_out = 8'h1E;
                    16'hB756: data_out = 8'h1F;
                    16'hB757: data_out = 8'h20;
                    16'hB758: data_out = 8'h21;
                    16'hB759: data_out = 8'h22;
                    16'hB75A: data_out = 8'h23;
                    16'hB75B: data_out = 8'h24;
                    16'hB75C: data_out = 8'h25;
                    16'hB75D: data_out = 8'h26;
                    16'hB75E: data_out = 8'h27;
                    16'hB75F: data_out = 8'h28;
                    16'hB760: data_out = 8'h29;
                    16'hB761: data_out = 8'h2A;
                    16'hB762: data_out = 8'h2B;
                    16'hB763: data_out = 8'h2C;
                    16'hB764: data_out = 8'h2D;
                    16'hB765: data_out = 8'h2E;
                    16'hB766: data_out = 8'h2F;
                    16'hB767: data_out = 8'h30;
                    16'hB768: data_out = 8'h31;
                    16'hB769: data_out = 8'h32;
                    16'hB76A: data_out = 8'h33;
                    16'hB76B: data_out = 8'h34;
                    16'hB76C: data_out = 8'h35;
                    16'hB76D: data_out = 8'h36;
                    16'hB76E: data_out = 8'h37;
                    16'hB76F: data_out = 8'h38;
                    16'hB770: data_out = 8'h39;
                    16'hB771: data_out = 8'h3A;
                    16'hB772: data_out = 8'h3B;
                    16'hB773: data_out = 8'h3C;
                    16'hB774: data_out = 8'h3D;
                    16'hB775: data_out = 8'h3E;
                    16'hB776: data_out = 8'h3F;
                    16'hB777: data_out = 8'h40;
                    16'hB778: data_out = 8'h41;
                    16'hB779: data_out = 8'h42;
                    16'hB77A: data_out = 8'h43;
                    16'hB77B: data_out = 8'h44;
                    16'hB77C: data_out = 8'h45;
                    16'hB77D: data_out = 8'h46;
                    16'hB77E: data_out = 8'h47;
                    16'hB77F: data_out = 8'h48;
                    16'hB780: data_out = 8'hB7;
                    16'hB781: data_out = 8'hB8;
                    16'hB782: data_out = 8'hB9;
                    16'hB783: data_out = 8'hBA;
                    16'hB784: data_out = 8'hBB;
                    16'hB785: data_out = 8'hBC;
                    16'hB786: data_out = 8'hBD;
                    16'hB787: data_out = 8'hBE;
                    16'hB788: data_out = 8'hBF;
                    16'hB789: data_out = 8'hC0;
                    16'hB78A: data_out = 8'hC1;
                    16'hB78B: data_out = 8'hC2;
                    16'hB78C: data_out = 8'hC3;
                    16'hB78D: data_out = 8'hC4;
                    16'hB78E: data_out = 8'hC5;
                    16'hB78F: data_out = 8'hC6;
                    16'hB790: data_out = 8'hC7;
                    16'hB791: data_out = 8'hC8;
                    16'hB792: data_out = 8'hC9;
                    16'hB793: data_out = 8'hCA;
                    16'hB794: data_out = 8'hCB;
                    16'hB795: data_out = 8'hCC;
                    16'hB796: data_out = 8'hCD;
                    16'hB797: data_out = 8'hCE;
                    16'hB798: data_out = 8'hCF;
                    16'hB799: data_out = 8'hD0;
                    16'hB79A: data_out = 8'hD1;
                    16'hB79B: data_out = 8'hD2;
                    16'hB79C: data_out = 8'hD3;
                    16'hB79D: data_out = 8'hD4;
                    16'hB79E: data_out = 8'hD5;
                    16'hB79F: data_out = 8'hD6;
                    16'hB7A0: data_out = 8'hD7;
                    16'hB7A1: data_out = 8'hD8;
                    16'hB7A2: data_out = 8'hD9;
                    16'hB7A3: data_out = 8'hDA;
                    16'hB7A4: data_out = 8'hDB;
                    16'hB7A5: data_out = 8'hDC;
                    16'hB7A6: data_out = 8'hDD;
                    16'hB7A7: data_out = 8'hDE;
                    16'hB7A8: data_out = 8'hDF;
                    16'hB7A9: data_out = 8'hE0;
                    16'hB7AA: data_out = 8'hE1;
                    16'hB7AB: data_out = 8'hE2;
                    16'hB7AC: data_out = 8'hE3;
                    16'hB7AD: data_out = 8'hE4;
                    16'hB7AE: data_out = 8'hE5;
                    16'hB7AF: data_out = 8'hE6;
                    16'hB7B0: data_out = 8'hE7;
                    16'hB7B1: data_out = 8'hE8;
                    16'hB7B2: data_out = 8'hE9;
                    16'hB7B3: data_out = 8'hEA;
                    16'hB7B4: data_out = 8'hEB;
                    16'hB7B5: data_out = 8'hEC;
                    16'hB7B6: data_out = 8'hED;
                    16'hB7B7: data_out = 8'hEE;
                    16'hB7B8: data_out = 8'hEF;
                    16'hB7B9: data_out = 8'hF0;
                    16'hB7BA: data_out = 8'hF1;
                    16'hB7BB: data_out = 8'hF2;
                    16'hB7BC: data_out = 8'hF3;
                    16'hB7BD: data_out = 8'hF4;
                    16'hB7BE: data_out = 8'hF5;
                    16'hB7BF: data_out = 8'hF6;
                    16'hB7C0: data_out = 8'hF7;
                    16'hB7C1: data_out = 8'hF8;
                    16'hB7C2: data_out = 8'hF9;
                    16'hB7C3: data_out = 8'hFA;
                    16'hB7C4: data_out = 8'hFB;
                    16'hB7C5: data_out = 8'hFC;
                    16'hB7C6: data_out = 8'hFD;
                    16'hB7C7: data_out = 8'hFE;
                    16'hB7C8: data_out = 8'hFF;
                    16'hB7C9: data_out = 8'h80;
                    16'hB7CA: data_out = 8'h81;
                    16'hB7CB: data_out = 8'h82;
                    16'hB7CC: data_out = 8'h83;
                    16'hB7CD: data_out = 8'h84;
                    16'hB7CE: data_out = 8'h85;
                    16'hB7CF: data_out = 8'h86;
                    16'hB7D0: data_out = 8'h87;
                    16'hB7D1: data_out = 8'h88;
                    16'hB7D2: data_out = 8'h89;
                    16'hB7D3: data_out = 8'h8A;
                    16'hB7D4: data_out = 8'h8B;
                    16'hB7D5: data_out = 8'h8C;
                    16'hB7D6: data_out = 8'h8D;
                    16'hB7D7: data_out = 8'h8E;
                    16'hB7D8: data_out = 8'h8F;
                    16'hB7D9: data_out = 8'h90;
                    16'hB7DA: data_out = 8'h91;
                    16'hB7DB: data_out = 8'h92;
                    16'hB7DC: data_out = 8'h93;
                    16'hB7DD: data_out = 8'h94;
                    16'hB7DE: data_out = 8'h95;
                    16'hB7DF: data_out = 8'h96;
                    16'hB7E0: data_out = 8'h97;
                    16'hB7E1: data_out = 8'h98;
                    16'hB7E2: data_out = 8'h99;
                    16'hB7E3: data_out = 8'h9A;
                    16'hB7E4: data_out = 8'h9B;
                    16'hB7E5: data_out = 8'h9C;
                    16'hB7E6: data_out = 8'h9D;
                    16'hB7E7: data_out = 8'h9E;
                    16'hB7E8: data_out = 8'h9F;
                    16'hB7E9: data_out = 8'hA0;
                    16'hB7EA: data_out = 8'hA1;
                    16'hB7EB: data_out = 8'hA2;
                    16'hB7EC: data_out = 8'hA3;
                    16'hB7ED: data_out = 8'hA4;
                    16'hB7EE: data_out = 8'hA5;
                    16'hB7EF: data_out = 8'hA6;
                    16'hB7F0: data_out = 8'hA7;
                    16'hB7F1: data_out = 8'hA8;
                    16'hB7F2: data_out = 8'hA9;
                    16'hB7F3: data_out = 8'hAA;
                    16'hB7F4: data_out = 8'hAB;
                    16'hB7F5: data_out = 8'hAC;
                    16'hB7F6: data_out = 8'hAD;
                    16'hB7F7: data_out = 8'hAE;
                    16'hB7F8: data_out = 8'hAF;
                    16'hB7F9: data_out = 8'hB0;
                    16'hB7FA: data_out = 8'hB1;
                    16'hB7FB: data_out = 8'hB2;
                    16'hB7FC: data_out = 8'hB3;
                    16'hB7FD: data_out = 8'hB4;
                    16'hB7FE: data_out = 8'hB5;
                    16'hB7FF: data_out = 8'hB6;
                    16'hB800: data_out = 8'hB8;
                    16'hB801: data_out = 8'hB7;
                    16'hB802: data_out = 8'hB6;
                    16'hB803: data_out = 8'hB5;
                    16'hB804: data_out = 8'hB4;
                    16'hB805: data_out = 8'hB3;
                    16'hB806: data_out = 8'hB2;
                    16'hB807: data_out = 8'hB1;
                    16'hB808: data_out = 8'hB0;
                    16'hB809: data_out = 8'hAF;
                    16'hB80A: data_out = 8'hAE;
                    16'hB80B: data_out = 8'hAD;
                    16'hB80C: data_out = 8'hAC;
                    16'hB80D: data_out = 8'hAB;
                    16'hB80E: data_out = 8'hAA;
                    16'hB80F: data_out = 8'hA9;
                    16'hB810: data_out = 8'hA8;
                    16'hB811: data_out = 8'hA7;
                    16'hB812: data_out = 8'hA6;
                    16'hB813: data_out = 8'hA5;
                    16'hB814: data_out = 8'hA4;
                    16'hB815: data_out = 8'hA3;
                    16'hB816: data_out = 8'hA2;
                    16'hB817: data_out = 8'hA1;
                    16'hB818: data_out = 8'hA0;
                    16'hB819: data_out = 8'h9F;
                    16'hB81A: data_out = 8'h9E;
                    16'hB81B: data_out = 8'h9D;
                    16'hB81C: data_out = 8'h9C;
                    16'hB81D: data_out = 8'h9B;
                    16'hB81E: data_out = 8'h9A;
                    16'hB81F: data_out = 8'h99;
                    16'hB820: data_out = 8'h98;
                    16'hB821: data_out = 8'h97;
                    16'hB822: data_out = 8'h96;
                    16'hB823: data_out = 8'h95;
                    16'hB824: data_out = 8'h94;
                    16'hB825: data_out = 8'h93;
                    16'hB826: data_out = 8'h92;
                    16'hB827: data_out = 8'h91;
                    16'hB828: data_out = 8'h90;
                    16'hB829: data_out = 8'h8F;
                    16'hB82A: data_out = 8'h8E;
                    16'hB82B: data_out = 8'h8D;
                    16'hB82C: data_out = 8'h8C;
                    16'hB82D: data_out = 8'h8B;
                    16'hB82E: data_out = 8'h8A;
                    16'hB82F: data_out = 8'h89;
                    16'hB830: data_out = 8'h88;
                    16'hB831: data_out = 8'h87;
                    16'hB832: data_out = 8'h86;
                    16'hB833: data_out = 8'h85;
                    16'hB834: data_out = 8'h84;
                    16'hB835: data_out = 8'h83;
                    16'hB836: data_out = 8'h82;
                    16'hB837: data_out = 8'h81;
                    16'hB838: data_out = 8'h0;
                    16'hB839: data_out = 8'h1;
                    16'hB83A: data_out = 8'h2;
                    16'hB83B: data_out = 8'h3;
                    16'hB83C: data_out = 8'h4;
                    16'hB83D: data_out = 8'h5;
                    16'hB83E: data_out = 8'h6;
                    16'hB83F: data_out = 8'h7;
                    16'hB840: data_out = 8'h8;
                    16'hB841: data_out = 8'h9;
                    16'hB842: data_out = 8'hA;
                    16'hB843: data_out = 8'hB;
                    16'hB844: data_out = 8'hC;
                    16'hB845: data_out = 8'hD;
                    16'hB846: data_out = 8'hE;
                    16'hB847: data_out = 8'hF;
                    16'hB848: data_out = 8'h10;
                    16'hB849: data_out = 8'h11;
                    16'hB84A: data_out = 8'h12;
                    16'hB84B: data_out = 8'h13;
                    16'hB84C: data_out = 8'h14;
                    16'hB84D: data_out = 8'h15;
                    16'hB84E: data_out = 8'h16;
                    16'hB84F: data_out = 8'h17;
                    16'hB850: data_out = 8'h18;
                    16'hB851: data_out = 8'h19;
                    16'hB852: data_out = 8'h1A;
                    16'hB853: data_out = 8'h1B;
                    16'hB854: data_out = 8'h1C;
                    16'hB855: data_out = 8'h1D;
                    16'hB856: data_out = 8'h1E;
                    16'hB857: data_out = 8'h1F;
                    16'hB858: data_out = 8'h20;
                    16'hB859: data_out = 8'h21;
                    16'hB85A: data_out = 8'h22;
                    16'hB85B: data_out = 8'h23;
                    16'hB85C: data_out = 8'h24;
                    16'hB85D: data_out = 8'h25;
                    16'hB85E: data_out = 8'h26;
                    16'hB85F: data_out = 8'h27;
                    16'hB860: data_out = 8'h28;
                    16'hB861: data_out = 8'h29;
                    16'hB862: data_out = 8'h2A;
                    16'hB863: data_out = 8'h2B;
                    16'hB864: data_out = 8'h2C;
                    16'hB865: data_out = 8'h2D;
                    16'hB866: data_out = 8'h2E;
                    16'hB867: data_out = 8'h2F;
                    16'hB868: data_out = 8'h30;
                    16'hB869: data_out = 8'h31;
                    16'hB86A: data_out = 8'h32;
                    16'hB86B: data_out = 8'h33;
                    16'hB86C: data_out = 8'h34;
                    16'hB86D: data_out = 8'h35;
                    16'hB86E: data_out = 8'h36;
                    16'hB86F: data_out = 8'h37;
                    16'hB870: data_out = 8'h38;
                    16'hB871: data_out = 8'h39;
                    16'hB872: data_out = 8'h3A;
                    16'hB873: data_out = 8'h3B;
                    16'hB874: data_out = 8'h3C;
                    16'hB875: data_out = 8'h3D;
                    16'hB876: data_out = 8'h3E;
                    16'hB877: data_out = 8'h3F;
                    16'hB878: data_out = 8'h40;
                    16'hB879: data_out = 8'h41;
                    16'hB87A: data_out = 8'h42;
                    16'hB87B: data_out = 8'h43;
                    16'hB87C: data_out = 8'h44;
                    16'hB87D: data_out = 8'h45;
                    16'hB87E: data_out = 8'h46;
                    16'hB87F: data_out = 8'h47;
                    16'hB880: data_out = 8'hB8;
                    16'hB881: data_out = 8'hB9;
                    16'hB882: data_out = 8'hBA;
                    16'hB883: data_out = 8'hBB;
                    16'hB884: data_out = 8'hBC;
                    16'hB885: data_out = 8'hBD;
                    16'hB886: data_out = 8'hBE;
                    16'hB887: data_out = 8'hBF;
                    16'hB888: data_out = 8'hC0;
                    16'hB889: data_out = 8'hC1;
                    16'hB88A: data_out = 8'hC2;
                    16'hB88B: data_out = 8'hC3;
                    16'hB88C: data_out = 8'hC4;
                    16'hB88D: data_out = 8'hC5;
                    16'hB88E: data_out = 8'hC6;
                    16'hB88F: data_out = 8'hC7;
                    16'hB890: data_out = 8'hC8;
                    16'hB891: data_out = 8'hC9;
                    16'hB892: data_out = 8'hCA;
                    16'hB893: data_out = 8'hCB;
                    16'hB894: data_out = 8'hCC;
                    16'hB895: data_out = 8'hCD;
                    16'hB896: data_out = 8'hCE;
                    16'hB897: data_out = 8'hCF;
                    16'hB898: data_out = 8'hD0;
                    16'hB899: data_out = 8'hD1;
                    16'hB89A: data_out = 8'hD2;
                    16'hB89B: data_out = 8'hD3;
                    16'hB89C: data_out = 8'hD4;
                    16'hB89D: data_out = 8'hD5;
                    16'hB89E: data_out = 8'hD6;
                    16'hB89F: data_out = 8'hD7;
                    16'hB8A0: data_out = 8'hD8;
                    16'hB8A1: data_out = 8'hD9;
                    16'hB8A2: data_out = 8'hDA;
                    16'hB8A3: data_out = 8'hDB;
                    16'hB8A4: data_out = 8'hDC;
                    16'hB8A5: data_out = 8'hDD;
                    16'hB8A6: data_out = 8'hDE;
                    16'hB8A7: data_out = 8'hDF;
                    16'hB8A8: data_out = 8'hE0;
                    16'hB8A9: data_out = 8'hE1;
                    16'hB8AA: data_out = 8'hE2;
                    16'hB8AB: data_out = 8'hE3;
                    16'hB8AC: data_out = 8'hE4;
                    16'hB8AD: data_out = 8'hE5;
                    16'hB8AE: data_out = 8'hE6;
                    16'hB8AF: data_out = 8'hE7;
                    16'hB8B0: data_out = 8'hE8;
                    16'hB8B1: data_out = 8'hE9;
                    16'hB8B2: data_out = 8'hEA;
                    16'hB8B3: data_out = 8'hEB;
                    16'hB8B4: data_out = 8'hEC;
                    16'hB8B5: data_out = 8'hED;
                    16'hB8B6: data_out = 8'hEE;
                    16'hB8B7: data_out = 8'hEF;
                    16'hB8B8: data_out = 8'hF0;
                    16'hB8B9: data_out = 8'hF1;
                    16'hB8BA: data_out = 8'hF2;
                    16'hB8BB: data_out = 8'hF3;
                    16'hB8BC: data_out = 8'hF4;
                    16'hB8BD: data_out = 8'hF5;
                    16'hB8BE: data_out = 8'hF6;
                    16'hB8BF: data_out = 8'hF7;
                    16'hB8C0: data_out = 8'hF8;
                    16'hB8C1: data_out = 8'hF9;
                    16'hB8C2: data_out = 8'hFA;
                    16'hB8C3: data_out = 8'hFB;
                    16'hB8C4: data_out = 8'hFC;
                    16'hB8C5: data_out = 8'hFD;
                    16'hB8C6: data_out = 8'hFE;
                    16'hB8C7: data_out = 8'hFF;
                    16'hB8C8: data_out = 8'h80;
                    16'hB8C9: data_out = 8'h81;
                    16'hB8CA: data_out = 8'h82;
                    16'hB8CB: data_out = 8'h83;
                    16'hB8CC: data_out = 8'h84;
                    16'hB8CD: data_out = 8'h85;
                    16'hB8CE: data_out = 8'h86;
                    16'hB8CF: data_out = 8'h87;
                    16'hB8D0: data_out = 8'h88;
                    16'hB8D1: data_out = 8'h89;
                    16'hB8D2: data_out = 8'h8A;
                    16'hB8D3: data_out = 8'h8B;
                    16'hB8D4: data_out = 8'h8C;
                    16'hB8D5: data_out = 8'h8D;
                    16'hB8D6: data_out = 8'h8E;
                    16'hB8D7: data_out = 8'h8F;
                    16'hB8D8: data_out = 8'h90;
                    16'hB8D9: data_out = 8'h91;
                    16'hB8DA: data_out = 8'h92;
                    16'hB8DB: data_out = 8'h93;
                    16'hB8DC: data_out = 8'h94;
                    16'hB8DD: data_out = 8'h95;
                    16'hB8DE: data_out = 8'h96;
                    16'hB8DF: data_out = 8'h97;
                    16'hB8E0: data_out = 8'h98;
                    16'hB8E1: data_out = 8'h99;
                    16'hB8E2: data_out = 8'h9A;
                    16'hB8E3: data_out = 8'h9B;
                    16'hB8E4: data_out = 8'h9C;
                    16'hB8E5: data_out = 8'h9D;
                    16'hB8E6: data_out = 8'h9E;
                    16'hB8E7: data_out = 8'h9F;
                    16'hB8E8: data_out = 8'hA0;
                    16'hB8E9: data_out = 8'hA1;
                    16'hB8EA: data_out = 8'hA2;
                    16'hB8EB: data_out = 8'hA3;
                    16'hB8EC: data_out = 8'hA4;
                    16'hB8ED: data_out = 8'hA5;
                    16'hB8EE: data_out = 8'hA6;
                    16'hB8EF: data_out = 8'hA7;
                    16'hB8F0: data_out = 8'hA8;
                    16'hB8F1: data_out = 8'hA9;
                    16'hB8F2: data_out = 8'hAA;
                    16'hB8F3: data_out = 8'hAB;
                    16'hB8F4: data_out = 8'hAC;
                    16'hB8F5: data_out = 8'hAD;
                    16'hB8F6: data_out = 8'hAE;
                    16'hB8F7: data_out = 8'hAF;
                    16'hB8F8: data_out = 8'hB0;
                    16'hB8F9: data_out = 8'hB1;
                    16'hB8FA: data_out = 8'hB2;
                    16'hB8FB: data_out = 8'hB3;
                    16'hB8FC: data_out = 8'hB4;
                    16'hB8FD: data_out = 8'hB5;
                    16'hB8FE: data_out = 8'hB6;
                    16'hB8FF: data_out = 8'hB7;
                    16'hB900: data_out = 8'hB9;
                    16'hB901: data_out = 8'hB8;
                    16'hB902: data_out = 8'hB7;
                    16'hB903: data_out = 8'hB6;
                    16'hB904: data_out = 8'hB5;
                    16'hB905: data_out = 8'hB4;
                    16'hB906: data_out = 8'hB3;
                    16'hB907: data_out = 8'hB2;
                    16'hB908: data_out = 8'hB1;
                    16'hB909: data_out = 8'hB0;
                    16'hB90A: data_out = 8'hAF;
                    16'hB90B: data_out = 8'hAE;
                    16'hB90C: data_out = 8'hAD;
                    16'hB90D: data_out = 8'hAC;
                    16'hB90E: data_out = 8'hAB;
                    16'hB90F: data_out = 8'hAA;
                    16'hB910: data_out = 8'hA9;
                    16'hB911: data_out = 8'hA8;
                    16'hB912: data_out = 8'hA7;
                    16'hB913: data_out = 8'hA6;
                    16'hB914: data_out = 8'hA5;
                    16'hB915: data_out = 8'hA4;
                    16'hB916: data_out = 8'hA3;
                    16'hB917: data_out = 8'hA2;
                    16'hB918: data_out = 8'hA1;
                    16'hB919: data_out = 8'hA0;
                    16'hB91A: data_out = 8'h9F;
                    16'hB91B: data_out = 8'h9E;
                    16'hB91C: data_out = 8'h9D;
                    16'hB91D: data_out = 8'h9C;
                    16'hB91E: data_out = 8'h9B;
                    16'hB91F: data_out = 8'h9A;
                    16'hB920: data_out = 8'h99;
                    16'hB921: data_out = 8'h98;
                    16'hB922: data_out = 8'h97;
                    16'hB923: data_out = 8'h96;
                    16'hB924: data_out = 8'h95;
                    16'hB925: data_out = 8'h94;
                    16'hB926: data_out = 8'h93;
                    16'hB927: data_out = 8'h92;
                    16'hB928: data_out = 8'h91;
                    16'hB929: data_out = 8'h90;
                    16'hB92A: data_out = 8'h8F;
                    16'hB92B: data_out = 8'h8E;
                    16'hB92C: data_out = 8'h8D;
                    16'hB92D: data_out = 8'h8C;
                    16'hB92E: data_out = 8'h8B;
                    16'hB92F: data_out = 8'h8A;
                    16'hB930: data_out = 8'h89;
                    16'hB931: data_out = 8'h88;
                    16'hB932: data_out = 8'h87;
                    16'hB933: data_out = 8'h86;
                    16'hB934: data_out = 8'h85;
                    16'hB935: data_out = 8'h84;
                    16'hB936: data_out = 8'h83;
                    16'hB937: data_out = 8'h82;
                    16'hB938: data_out = 8'h81;
                    16'hB939: data_out = 8'h0;
                    16'hB93A: data_out = 8'h1;
                    16'hB93B: data_out = 8'h2;
                    16'hB93C: data_out = 8'h3;
                    16'hB93D: data_out = 8'h4;
                    16'hB93E: data_out = 8'h5;
                    16'hB93F: data_out = 8'h6;
                    16'hB940: data_out = 8'h7;
                    16'hB941: data_out = 8'h8;
                    16'hB942: data_out = 8'h9;
                    16'hB943: data_out = 8'hA;
                    16'hB944: data_out = 8'hB;
                    16'hB945: data_out = 8'hC;
                    16'hB946: data_out = 8'hD;
                    16'hB947: data_out = 8'hE;
                    16'hB948: data_out = 8'hF;
                    16'hB949: data_out = 8'h10;
                    16'hB94A: data_out = 8'h11;
                    16'hB94B: data_out = 8'h12;
                    16'hB94C: data_out = 8'h13;
                    16'hB94D: data_out = 8'h14;
                    16'hB94E: data_out = 8'h15;
                    16'hB94F: data_out = 8'h16;
                    16'hB950: data_out = 8'h17;
                    16'hB951: data_out = 8'h18;
                    16'hB952: data_out = 8'h19;
                    16'hB953: data_out = 8'h1A;
                    16'hB954: data_out = 8'h1B;
                    16'hB955: data_out = 8'h1C;
                    16'hB956: data_out = 8'h1D;
                    16'hB957: data_out = 8'h1E;
                    16'hB958: data_out = 8'h1F;
                    16'hB959: data_out = 8'h20;
                    16'hB95A: data_out = 8'h21;
                    16'hB95B: data_out = 8'h22;
                    16'hB95C: data_out = 8'h23;
                    16'hB95D: data_out = 8'h24;
                    16'hB95E: data_out = 8'h25;
                    16'hB95F: data_out = 8'h26;
                    16'hB960: data_out = 8'h27;
                    16'hB961: data_out = 8'h28;
                    16'hB962: data_out = 8'h29;
                    16'hB963: data_out = 8'h2A;
                    16'hB964: data_out = 8'h2B;
                    16'hB965: data_out = 8'h2C;
                    16'hB966: data_out = 8'h2D;
                    16'hB967: data_out = 8'h2E;
                    16'hB968: data_out = 8'h2F;
                    16'hB969: data_out = 8'h30;
                    16'hB96A: data_out = 8'h31;
                    16'hB96B: data_out = 8'h32;
                    16'hB96C: data_out = 8'h33;
                    16'hB96D: data_out = 8'h34;
                    16'hB96E: data_out = 8'h35;
                    16'hB96F: data_out = 8'h36;
                    16'hB970: data_out = 8'h37;
                    16'hB971: data_out = 8'h38;
                    16'hB972: data_out = 8'h39;
                    16'hB973: data_out = 8'h3A;
                    16'hB974: data_out = 8'h3B;
                    16'hB975: data_out = 8'h3C;
                    16'hB976: data_out = 8'h3D;
                    16'hB977: data_out = 8'h3E;
                    16'hB978: data_out = 8'h3F;
                    16'hB979: data_out = 8'h40;
                    16'hB97A: data_out = 8'h41;
                    16'hB97B: data_out = 8'h42;
                    16'hB97C: data_out = 8'h43;
                    16'hB97D: data_out = 8'h44;
                    16'hB97E: data_out = 8'h45;
                    16'hB97F: data_out = 8'h46;
                    16'hB980: data_out = 8'hB9;
                    16'hB981: data_out = 8'hBA;
                    16'hB982: data_out = 8'hBB;
                    16'hB983: data_out = 8'hBC;
                    16'hB984: data_out = 8'hBD;
                    16'hB985: data_out = 8'hBE;
                    16'hB986: data_out = 8'hBF;
                    16'hB987: data_out = 8'hC0;
                    16'hB988: data_out = 8'hC1;
                    16'hB989: data_out = 8'hC2;
                    16'hB98A: data_out = 8'hC3;
                    16'hB98B: data_out = 8'hC4;
                    16'hB98C: data_out = 8'hC5;
                    16'hB98D: data_out = 8'hC6;
                    16'hB98E: data_out = 8'hC7;
                    16'hB98F: data_out = 8'hC8;
                    16'hB990: data_out = 8'hC9;
                    16'hB991: data_out = 8'hCA;
                    16'hB992: data_out = 8'hCB;
                    16'hB993: data_out = 8'hCC;
                    16'hB994: data_out = 8'hCD;
                    16'hB995: data_out = 8'hCE;
                    16'hB996: data_out = 8'hCF;
                    16'hB997: data_out = 8'hD0;
                    16'hB998: data_out = 8'hD1;
                    16'hB999: data_out = 8'hD2;
                    16'hB99A: data_out = 8'hD3;
                    16'hB99B: data_out = 8'hD4;
                    16'hB99C: data_out = 8'hD5;
                    16'hB99D: data_out = 8'hD6;
                    16'hB99E: data_out = 8'hD7;
                    16'hB99F: data_out = 8'hD8;
                    16'hB9A0: data_out = 8'hD9;
                    16'hB9A1: data_out = 8'hDA;
                    16'hB9A2: data_out = 8'hDB;
                    16'hB9A3: data_out = 8'hDC;
                    16'hB9A4: data_out = 8'hDD;
                    16'hB9A5: data_out = 8'hDE;
                    16'hB9A6: data_out = 8'hDF;
                    16'hB9A7: data_out = 8'hE0;
                    16'hB9A8: data_out = 8'hE1;
                    16'hB9A9: data_out = 8'hE2;
                    16'hB9AA: data_out = 8'hE3;
                    16'hB9AB: data_out = 8'hE4;
                    16'hB9AC: data_out = 8'hE5;
                    16'hB9AD: data_out = 8'hE6;
                    16'hB9AE: data_out = 8'hE7;
                    16'hB9AF: data_out = 8'hE8;
                    16'hB9B0: data_out = 8'hE9;
                    16'hB9B1: data_out = 8'hEA;
                    16'hB9B2: data_out = 8'hEB;
                    16'hB9B3: data_out = 8'hEC;
                    16'hB9B4: data_out = 8'hED;
                    16'hB9B5: data_out = 8'hEE;
                    16'hB9B6: data_out = 8'hEF;
                    16'hB9B7: data_out = 8'hF0;
                    16'hB9B8: data_out = 8'hF1;
                    16'hB9B9: data_out = 8'hF2;
                    16'hB9BA: data_out = 8'hF3;
                    16'hB9BB: data_out = 8'hF4;
                    16'hB9BC: data_out = 8'hF5;
                    16'hB9BD: data_out = 8'hF6;
                    16'hB9BE: data_out = 8'hF7;
                    16'hB9BF: data_out = 8'hF8;
                    16'hB9C0: data_out = 8'hF9;
                    16'hB9C1: data_out = 8'hFA;
                    16'hB9C2: data_out = 8'hFB;
                    16'hB9C3: data_out = 8'hFC;
                    16'hB9C4: data_out = 8'hFD;
                    16'hB9C5: data_out = 8'hFE;
                    16'hB9C6: data_out = 8'hFF;
                    16'hB9C7: data_out = 8'h80;
                    16'hB9C8: data_out = 8'h81;
                    16'hB9C9: data_out = 8'h82;
                    16'hB9CA: data_out = 8'h83;
                    16'hB9CB: data_out = 8'h84;
                    16'hB9CC: data_out = 8'h85;
                    16'hB9CD: data_out = 8'h86;
                    16'hB9CE: data_out = 8'h87;
                    16'hB9CF: data_out = 8'h88;
                    16'hB9D0: data_out = 8'h89;
                    16'hB9D1: data_out = 8'h8A;
                    16'hB9D2: data_out = 8'h8B;
                    16'hB9D3: data_out = 8'h8C;
                    16'hB9D4: data_out = 8'h8D;
                    16'hB9D5: data_out = 8'h8E;
                    16'hB9D6: data_out = 8'h8F;
                    16'hB9D7: data_out = 8'h90;
                    16'hB9D8: data_out = 8'h91;
                    16'hB9D9: data_out = 8'h92;
                    16'hB9DA: data_out = 8'h93;
                    16'hB9DB: data_out = 8'h94;
                    16'hB9DC: data_out = 8'h95;
                    16'hB9DD: data_out = 8'h96;
                    16'hB9DE: data_out = 8'h97;
                    16'hB9DF: data_out = 8'h98;
                    16'hB9E0: data_out = 8'h99;
                    16'hB9E1: data_out = 8'h9A;
                    16'hB9E2: data_out = 8'h9B;
                    16'hB9E3: data_out = 8'h9C;
                    16'hB9E4: data_out = 8'h9D;
                    16'hB9E5: data_out = 8'h9E;
                    16'hB9E6: data_out = 8'h9F;
                    16'hB9E7: data_out = 8'hA0;
                    16'hB9E8: data_out = 8'hA1;
                    16'hB9E9: data_out = 8'hA2;
                    16'hB9EA: data_out = 8'hA3;
                    16'hB9EB: data_out = 8'hA4;
                    16'hB9EC: data_out = 8'hA5;
                    16'hB9ED: data_out = 8'hA6;
                    16'hB9EE: data_out = 8'hA7;
                    16'hB9EF: data_out = 8'hA8;
                    16'hB9F0: data_out = 8'hA9;
                    16'hB9F1: data_out = 8'hAA;
                    16'hB9F2: data_out = 8'hAB;
                    16'hB9F3: data_out = 8'hAC;
                    16'hB9F4: data_out = 8'hAD;
                    16'hB9F5: data_out = 8'hAE;
                    16'hB9F6: data_out = 8'hAF;
                    16'hB9F7: data_out = 8'hB0;
                    16'hB9F8: data_out = 8'hB1;
                    16'hB9F9: data_out = 8'hB2;
                    16'hB9FA: data_out = 8'hB3;
                    16'hB9FB: data_out = 8'hB4;
                    16'hB9FC: data_out = 8'hB5;
                    16'hB9FD: data_out = 8'hB6;
                    16'hB9FE: data_out = 8'hB7;
                    16'hB9FF: data_out = 8'hB8;
                    16'hBA00: data_out = 8'hBA;
                    16'hBA01: data_out = 8'hB9;
                    16'hBA02: data_out = 8'hB8;
                    16'hBA03: data_out = 8'hB7;
                    16'hBA04: data_out = 8'hB6;
                    16'hBA05: data_out = 8'hB5;
                    16'hBA06: data_out = 8'hB4;
                    16'hBA07: data_out = 8'hB3;
                    16'hBA08: data_out = 8'hB2;
                    16'hBA09: data_out = 8'hB1;
                    16'hBA0A: data_out = 8'hB0;
                    16'hBA0B: data_out = 8'hAF;
                    16'hBA0C: data_out = 8'hAE;
                    16'hBA0D: data_out = 8'hAD;
                    16'hBA0E: data_out = 8'hAC;
                    16'hBA0F: data_out = 8'hAB;
                    16'hBA10: data_out = 8'hAA;
                    16'hBA11: data_out = 8'hA9;
                    16'hBA12: data_out = 8'hA8;
                    16'hBA13: data_out = 8'hA7;
                    16'hBA14: data_out = 8'hA6;
                    16'hBA15: data_out = 8'hA5;
                    16'hBA16: data_out = 8'hA4;
                    16'hBA17: data_out = 8'hA3;
                    16'hBA18: data_out = 8'hA2;
                    16'hBA19: data_out = 8'hA1;
                    16'hBA1A: data_out = 8'hA0;
                    16'hBA1B: data_out = 8'h9F;
                    16'hBA1C: data_out = 8'h9E;
                    16'hBA1D: data_out = 8'h9D;
                    16'hBA1E: data_out = 8'h9C;
                    16'hBA1F: data_out = 8'h9B;
                    16'hBA20: data_out = 8'h9A;
                    16'hBA21: data_out = 8'h99;
                    16'hBA22: data_out = 8'h98;
                    16'hBA23: data_out = 8'h97;
                    16'hBA24: data_out = 8'h96;
                    16'hBA25: data_out = 8'h95;
                    16'hBA26: data_out = 8'h94;
                    16'hBA27: data_out = 8'h93;
                    16'hBA28: data_out = 8'h92;
                    16'hBA29: data_out = 8'h91;
                    16'hBA2A: data_out = 8'h90;
                    16'hBA2B: data_out = 8'h8F;
                    16'hBA2C: data_out = 8'h8E;
                    16'hBA2D: data_out = 8'h8D;
                    16'hBA2E: data_out = 8'h8C;
                    16'hBA2F: data_out = 8'h8B;
                    16'hBA30: data_out = 8'h8A;
                    16'hBA31: data_out = 8'h89;
                    16'hBA32: data_out = 8'h88;
                    16'hBA33: data_out = 8'h87;
                    16'hBA34: data_out = 8'h86;
                    16'hBA35: data_out = 8'h85;
                    16'hBA36: data_out = 8'h84;
                    16'hBA37: data_out = 8'h83;
                    16'hBA38: data_out = 8'h82;
                    16'hBA39: data_out = 8'h81;
                    16'hBA3A: data_out = 8'h0;
                    16'hBA3B: data_out = 8'h1;
                    16'hBA3C: data_out = 8'h2;
                    16'hBA3D: data_out = 8'h3;
                    16'hBA3E: data_out = 8'h4;
                    16'hBA3F: data_out = 8'h5;
                    16'hBA40: data_out = 8'h6;
                    16'hBA41: data_out = 8'h7;
                    16'hBA42: data_out = 8'h8;
                    16'hBA43: data_out = 8'h9;
                    16'hBA44: data_out = 8'hA;
                    16'hBA45: data_out = 8'hB;
                    16'hBA46: data_out = 8'hC;
                    16'hBA47: data_out = 8'hD;
                    16'hBA48: data_out = 8'hE;
                    16'hBA49: data_out = 8'hF;
                    16'hBA4A: data_out = 8'h10;
                    16'hBA4B: data_out = 8'h11;
                    16'hBA4C: data_out = 8'h12;
                    16'hBA4D: data_out = 8'h13;
                    16'hBA4E: data_out = 8'h14;
                    16'hBA4F: data_out = 8'h15;
                    16'hBA50: data_out = 8'h16;
                    16'hBA51: data_out = 8'h17;
                    16'hBA52: data_out = 8'h18;
                    16'hBA53: data_out = 8'h19;
                    16'hBA54: data_out = 8'h1A;
                    16'hBA55: data_out = 8'h1B;
                    16'hBA56: data_out = 8'h1C;
                    16'hBA57: data_out = 8'h1D;
                    16'hBA58: data_out = 8'h1E;
                    16'hBA59: data_out = 8'h1F;
                    16'hBA5A: data_out = 8'h20;
                    16'hBA5B: data_out = 8'h21;
                    16'hBA5C: data_out = 8'h22;
                    16'hBA5D: data_out = 8'h23;
                    16'hBA5E: data_out = 8'h24;
                    16'hBA5F: data_out = 8'h25;
                    16'hBA60: data_out = 8'h26;
                    16'hBA61: data_out = 8'h27;
                    16'hBA62: data_out = 8'h28;
                    16'hBA63: data_out = 8'h29;
                    16'hBA64: data_out = 8'h2A;
                    16'hBA65: data_out = 8'h2B;
                    16'hBA66: data_out = 8'h2C;
                    16'hBA67: data_out = 8'h2D;
                    16'hBA68: data_out = 8'h2E;
                    16'hBA69: data_out = 8'h2F;
                    16'hBA6A: data_out = 8'h30;
                    16'hBA6B: data_out = 8'h31;
                    16'hBA6C: data_out = 8'h32;
                    16'hBA6D: data_out = 8'h33;
                    16'hBA6E: data_out = 8'h34;
                    16'hBA6F: data_out = 8'h35;
                    16'hBA70: data_out = 8'h36;
                    16'hBA71: data_out = 8'h37;
                    16'hBA72: data_out = 8'h38;
                    16'hBA73: data_out = 8'h39;
                    16'hBA74: data_out = 8'h3A;
                    16'hBA75: data_out = 8'h3B;
                    16'hBA76: data_out = 8'h3C;
                    16'hBA77: data_out = 8'h3D;
                    16'hBA78: data_out = 8'h3E;
                    16'hBA79: data_out = 8'h3F;
                    16'hBA7A: data_out = 8'h40;
                    16'hBA7B: data_out = 8'h41;
                    16'hBA7C: data_out = 8'h42;
                    16'hBA7D: data_out = 8'h43;
                    16'hBA7E: data_out = 8'h44;
                    16'hBA7F: data_out = 8'h45;
                    16'hBA80: data_out = 8'hBA;
                    16'hBA81: data_out = 8'hBB;
                    16'hBA82: data_out = 8'hBC;
                    16'hBA83: data_out = 8'hBD;
                    16'hBA84: data_out = 8'hBE;
                    16'hBA85: data_out = 8'hBF;
                    16'hBA86: data_out = 8'hC0;
                    16'hBA87: data_out = 8'hC1;
                    16'hBA88: data_out = 8'hC2;
                    16'hBA89: data_out = 8'hC3;
                    16'hBA8A: data_out = 8'hC4;
                    16'hBA8B: data_out = 8'hC5;
                    16'hBA8C: data_out = 8'hC6;
                    16'hBA8D: data_out = 8'hC7;
                    16'hBA8E: data_out = 8'hC8;
                    16'hBA8F: data_out = 8'hC9;
                    16'hBA90: data_out = 8'hCA;
                    16'hBA91: data_out = 8'hCB;
                    16'hBA92: data_out = 8'hCC;
                    16'hBA93: data_out = 8'hCD;
                    16'hBA94: data_out = 8'hCE;
                    16'hBA95: data_out = 8'hCF;
                    16'hBA96: data_out = 8'hD0;
                    16'hBA97: data_out = 8'hD1;
                    16'hBA98: data_out = 8'hD2;
                    16'hBA99: data_out = 8'hD3;
                    16'hBA9A: data_out = 8'hD4;
                    16'hBA9B: data_out = 8'hD5;
                    16'hBA9C: data_out = 8'hD6;
                    16'hBA9D: data_out = 8'hD7;
                    16'hBA9E: data_out = 8'hD8;
                    16'hBA9F: data_out = 8'hD9;
                    16'hBAA0: data_out = 8'hDA;
                    16'hBAA1: data_out = 8'hDB;
                    16'hBAA2: data_out = 8'hDC;
                    16'hBAA3: data_out = 8'hDD;
                    16'hBAA4: data_out = 8'hDE;
                    16'hBAA5: data_out = 8'hDF;
                    16'hBAA6: data_out = 8'hE0;
                    16'hBAA7: data_out = 8'hE1;
                    16'hBAA8: data_out = 8'hE2;
                    16'hBAA9: data_out = 8'hE3;
                    16'hBAAA: data_out = 8'hE4;
                    16'hBAAB: data_out = 8'hE5;
                    16'hBAAC: data_out = 8'hE6;
                    16'hBAAD: data_out = 8'hE7;
                    16'hBAAE: data_out = 8'hE8;
                    16'hBAAF: data_out = 8'hE9;
                    16'hBAB0: data_out = 8'hEA;
                    16'hBAB1: data_out = 8'hEB;
                    16'hBAB2: data_out = 8'hEC;
                    16'hBAB3: data_out = 8'hED;
                    16'hBAB4: data_out = 8'hEE;
                    16'hBAB5: data_out = 8'hEF;
                    16'hBAB6: data_out = 8'hF0;
                    16'hBAB7: data_out = 8'hF1;
                    16'hBAB8: data_out = 8'hF2;
                    16'hBAB9: data_out = 8'hF3;
                    16'hBABA: data_out = 8'hF4;
                    16'hBABB: data_out = 8'hF5;
                    16'hBABC: data_out = 8'hF6;
                    16'hBABD: data_out = 8'hF7;
                    16'hBABE: data_out = 8'hF8;
                    16'hBABF: data_out = 8'hF9;
                    16'hBAC0: data_out = 8'hFA;
                    16'hBAC1: data_out = 8'hFB;
                    16'hBAC2: data_out = 8'hFC;
                    16'hBAC3: data_out = 8'hFD;
                    16'hBAC4: data_out = 8'hFE;
                    16'hBAC5: data_out = 8'hFF;
                    16'hBAC6: data_out = 8'h80;
                    16'hBAC7: data_out = 8'h81;
                    16'hBAC8: data_out = 8'h82;
                    16'hBAC9: data_out = 8'h83;
                    16'hBACA: data_out = 8'h84;
                    16'hBACB: data_out = 8'h85;
                    16'hBACC: data_out = 8'h86;
                    16'hBACD: data_out = 8'h87;
                    16'hBACE: data_out = 8'h88;
                    16'hBACF: data_out = 8'h89;
                    16'hBAD0: data_out = 8'h8A;
                    16'hBAD1: data_out = 8'h8B;
                    16'hBAD2: data_out = 8'h8C;
                    16'hBAD3: data_out = 8'h8D;
                    16'hBAD4: data_out = 8'h8E;
                    16'hBAD5: data_out = 8'h8F;
                    16'hBAD6: data_out = 8'h90;
                    16'hBAD7: data_out = 8'h91;
                    16'hBAD8: data_out = 8'h92;
                    16'hBAD9: data_out = 8'h93;
                    16'hBADA: data_out = 8'h94;
                    16'hBADB: data_out = 8'h95;
                    16'hBADC: data_out = 8'h96;
                    16'hBADD: data_out = 8'h97;
                    16'hBADE: data_out = 8'h98;
                    16'hBADF: data_out = 8'h99;
                    16'hBAE0: data_out = 8'h9A;
                    16'hBAE1: data_out = 8'h9B;
                    16'hBAE2: data_out = 8'h9C;
                    16'hBAE3: data_out = 8'h9D;
                    16'hBAE4: data_out = 8'h9E;
                    16'hBAE5: data_out = 8'h9F;
                    16'hBAE6: data_out = 8'hA0;
                    16'hBAE7: data_out = 8'hA1;
                    16'hBAE8: data_out = 8'hA2;
                    16'hBAE9: data_out = 8'hA3;
                    16'hBAEA: data_out = 8'hA4;
                    16'hBAEB: data_out = 8'hA5;
                    16'hBAEC: data_out = 8'hA6;
                    16'hBAED: data_out = 8'hA7;
                    16'hBAEE: data_out = 8'hA8;
                    16'hBAEF: data_out = 8'hA9;
                    16'hBAF0: data_out = 8'hAA;
                    16'hBAF1: data_out = 8'hAB;
                    16'hBAF2: data_out = 8'hAC;
                    16'hBAF3: data_out = 8'hAD;
                    16'hBAF4: data_out = 8'hAE;
                    16'hBAF5: data_out = 8'hAF;
                    16'hBAF6: data_out = 8'hB0;
                    16'hBAF7: data_out = 8'hB1;
                    16'hBAF8: data_out = 8'hB2;
                    16'hBAF9: data_out = 8'hB3;
                    16'hBAFA: data_out = 8'hB4;
                    16'hBAFB: data_out = 8'hB5;
                    16'hBAFC: data_out = 8'hB6;
                    16'hBAFD: data_out = 8'hB7;
                    16'hBAFE: data_out = 8'hB8;
                    16'hBAFF: data_out = 8'hB9;
                    16'hBB00: data_out = 8'hBB;
                    16'hBB01: data_out = 8'hBA;
                    16'hBB02: data_out = 8'hB9;
                    16'hBB03: data_out = 8'hB8;
                    16'hBB04: data_out = 8'hB7;
                    16'hBB05: data_out = 8'hB6;
                    16'hBB06: data_out = 8'hB5;
                    16'hBB07: data_out = 8'hB4;
                    16'hBB08: data_out = 8'hB3;
                    16'hBB09: data_out = 8'hB2;
                    16'hBB0A: data_out = 8'hB1;
                    16'hBB0B: data_out = 8'hB0;
                    16'hBB0C: data_out = 8'hAF;
                    16'hBB0D: data_out = 8'hAE;
                    16'hBB0E: data_out = 8'hAD;
                    16'hBB0F: data_out = 8'hAC;
                    16'hBB10: data_out = 8'hAB;
                    16'hBB11: data_out = 8'hAA;
                    16'hBB12: data_out = 8'hA9;
                    16'hBB13: data_out = 8'hA8;
                    16'hBB14: data_out = 8'hA7;
                    16'hBB15: data_out = 8'hA6;
                    16'hBB16: data_out = 8'hA5;
                    16'hBB17: data_out = 8'hA4;
                    16'hBB18: data_out = 8'hA3;
                    16'hBB19: data_out = 8'hA2;
                    16'hBB1A: data_out = 8'hA1;
                    16'hBB1B: data_out = 8'hA0;
                    16'hBB1C: data_out = 8'h9F;
                    16'hBB1D: data_out = 8'h9E;
                    16'hBB1E: data_out = 8'h9D;
                    16'hBB1F: data_out = 8'h9C;
                    16'hBB20: data_out = 8'h9B;
                    16'hBB21: data_out = 8'h9A;
                    16'hBB22: data_out = 8'h99;
                    16'hBB23: data_out = 8'h98;
                    16'hBB24: data_out = 8'h97;
                    16'hBB25: data_out = 8'h96;
                    16'hBB26: data_out = 8'h95;
                    16'hBB27: data_out = 8'h94;
                    16'hBB28: data_out = 8'h93;
                    16'hBB29: data_out = 8'h92;
                    16'hBB2A: data_out = 8'h91;
                    16'hBB2B: data_out = 8'h90;
                    16'hBB2C: data_out = 8'h8F;
                    16'hBB2D: data_out = 8'h8E;
                    16'hBB2E: data_out = 8'h8D;
                    16'hBB2F: data_out = 8'h8C;
                    16'hBB30: data_out = 8'h8B;
                    16'hBB31: data_out = 8'h8A;
                    16'hBB32: data_out = 8'h89;
                    16'hBB33: data_out = 8'h88;
                    16'hBB34: data_out = 8'h87;
                    16'hBB35: data_out = 8'h86;
                    16'hBB36: data_out = 8'h85;
                    16'hBB37: data_out = 8'h84;
                    16'hBB38: data_out = 8'h83;
                    16'hBB39: data_out = 8'h82;
                    16'hBB3A: data_out = 8'h81;
                    16'hBB3B: data_out = 8'h0;
                    16'hBB3C: data_out = 8'h1;
                    16'hBB3D: data_out = 8'h2;
                    16'hBB3E: data_out = 8'h3;
                    16'hBB3F: data_out = 8'h4;
                    16'hBB40: data_out = 8'h5;
                    16'hBB41: data_out = 8'h6;
                    16'hBB42: data_out = 8'h7;
                    16'hBB43: data_out = 8'h8;
                    16'hBB44: data_out = 8'h9;
                    16'hBB45: data_out = 8'hA;
                    16'hBB46: data_out = 8'hB;
                    16'hBB47: data_out = 8'hC;
                    16'hBB48: data_out = 8'hD;
                    16'hBB49: data_out = 8'hE;
                    16'hBB4A: data_out = 8'hF;
                    16'hBB4B: data_out = 8'h10;
                    16'hBB4C: data_out = 8'h11;
                    16'hBB4D: data_out = 8'h12;
                    16'hBB4E: data_out = 8'h13;
                    16'hBB4F: data_out = 8'h14;
                    16'hBB50: data_out = 8'h15;
                    16'hBB51: data_out = 8'h16;
                    16'hBB52: data_out = 8'h17;
                    16'hBB53: data_out = 8'h18;
                    16'hBB54: data_out = 8'h19;
                    16'hBB55: data_out = 8'h1A;
                    16'hBB56: data_out = 8'h1B;
                    16'hBB57: data_out = 8'h1C;
                    16'hBB58: data_out = 8'h1D;
                    16'hBB59: data_out = 8'h1E;
                    16'hBB5A: data_out = 8'h1F;
                    16'hBB5B: data_out = 8'h20;
                    16'hBB5C: data_out = 8'h21;
                    16'hBB5D: data_out = 8'h22;
                    16'hBB5E: data_out = 8'h23;
                    16'hBB5F: data_out = 8'h24;
                    16'hBB60: data_out = 8'h25;
                    16'hBB61: data_out = 8'h26;
                    16'hBB62: data_out = 8'h27;
                    16'hBB63: data_out = 8'h28;
                    16'hBB64: data_out = 8'h29;
                    16'hBB65: data_out = 8'h2A;
                    16'hBB66: data_out = 8'h2B;
                    16'hBB67: data_out = 8'h2C;
                    16'hBB68: data_out = 8'h2D;
                    16'hBB69: data_out = 8'h2E;
                    16'hBB6A: data_out = 8'h2F;
                    16'hBB6B: data_out = 8'h30;
                    16'hBB6C: data_out = 8'h31;
                    16'hBB6D: data_out = 8'h32;
                    16'hBB6E: data_out = 8'h33;
                    16'hBB6F: data_out = 8'h34;
                    16'hBB70: data_out = 8'h35;
                    16'hBB71: data_out = 8'h36;
                    16'hBB72: data_out = 8'h37;
                    16'hBB73: data_out = 8'h38;
                    16'hBB74: data_out = 8'h39;
                    16'hBB75: data_out = 8'h3A;
                    16'hBB76: data_out = 8'h3B;
                    16'hBB77: data_out = 8'h3C;
                    16'hBB78: data_out = 8'h3D;
                    16'hBB79: data_out = 8'h3E;
                    16'hBB7A: data_out = 8'h3F;
                    16'hBB7B: data_out = 8'h40;
                    16'hBB7C: data_out = 8'h41;
                    16'hBB7D: data_out = 8'h42;
                    16'hBB7E: data_out = 8'h43;
                    16'hBB7F: data_out = 8'h44;
                    16'hBB80: data_out = 8'hBB;
                    16'hBB81: data_out = 8'hBC;
                    16'hBB82: data_out = 8'hBD;
                    16'hBB83: data_out = 8'hBE;
                    16'hBB84: data_out = 8'hBF;
                    16'hBB85: data_out = 8'hC0;
                    16'hBB86: data_out = 8'hC1;
                    16'hBB87: data_out = 8'hC2;
                    16'hBB88: data_out = 8'hC3;
                    16'hBB89: data_out = 8'hC4;
                    16'hBB8A: data_out = 8'hC5;
                    16'hBB8B: data_out = 8'hC6;
                    16'hBB8C: data_out = 8'hC7;
                    16'hBB8D: data_out = 8'hC8;
                    16'hBB8E: data_out = 8'hC9;
                    16'hBB8F: data_out = 8'hCA;
                    16'hBB90: data_out = 8'hCB;
                    16'hBB91: data_out = 8'hCC;
                    16'hBB92: data_out = 8'hCD;
                    16'hBB93: data_out = 8'hCE;
                    16'hBB94: data_out = 8'hCF;
                    16'hBB95: data_out = 8'hD0;
                    16'hBB96: data_out = 8'hD1;
                    16'hBB97: data_out = 8'hD2;
                    16'hBB98: data_out = 8'hD3;
                    16'hBB99: data_out = 8'hD4;
                    16'hBB9A: data_out = 8'hD5;
                    16'hBB9B: data_out = 8'hD6;
                    16'hBB9C: data_out = 8'hD7;
                    16'hBB9D: data_out = 8'hD8;
                    16'hBB9E: data_out = 8'hD9;
                    16'hBB9F: data_out = 8'hDA;
                    16'hBBA0: data_out = 8'hDB;
                    16'hBBA1: data_out = 8'hDC;
                    16'hBBA2: data_out = 8'hDD;
                    16'hBBA3: data_out = 8'hDE;
                    16'hBBA4: data_out = 8'hDF;
                    16'hBBA5: data_out = 8'hE0;
                    16'hBBA6: data_out = 8'hE1;
                    16'hBBA7: data_out = 8'hE2;
                    16'hBBA8: data_out = 8'hE3;
                    16'hBBA9: data_out = 8'hE4;
                    16'hBBAA: data_out = 8'hE5;
                    16'hBBAB: data_out = 8'hE6;
                    16'hBBAC: data_out = 8'hE7;
                    16'hBBAD: data_out = 8'hE8;
                    16'hBBAE: data_out = 8'hE9;
                    16'hBBAF: data_out = 8'hEA;
                    16'hBBB0: data_out = 8'hEB;
                    16'hBBB1: data_out = 8'hEC;
                    16'hBBB2: data_out = 8'hED;
                    16'hBBB3: data_out = 8'hEE;
                    16'hBBB4: data_out = 8'hEF;
                    16'hBBB5: data_out = 8'hF0;
                    16'hBBB6: data_out = 8'hF1;
                    16'hBBB7: data_out = 8'hF2;
                    16'hBBB8: data_out = 8'hF3;
                    16'hBBB9: data_out = 8'hF4;
                    16'hBBBA: data_out = 8'hF5;
                    16'hBBBB: data_out = 8'hF6;
                    16'hBBBC: data_out = 8'hF7;
                    16'hBBBD: data_out = 8'hF8;
                    16'hBBBE: data_out = 8'hF9;
                    16'hBBBF: data_out = 8'hFA;
                    16'hBBC0: data_out = 8'hFB;
                    16'hBBC1: data_out = 8'hFC;
                    16'hBBC2: data_out = 8'hFD;
                    16'hBBC3: data_out = 8'hFE;
                    16'hBBC4: data_out = 8'hFF;
                    16'hBBC5: data_out = 8'h80;
                    16'hBBC6: data_out = 8'h81;
                    16'hBBC7: data_out = 8'h82;
                    16'hBBC8: data_out = 8'h83;
                    16'hBBC9: data_out = 8'h84;
                    16'hBBCA: data_out = 8'h85;
                    16'hBBCB: data_out = 8'h86;
                    16'hBBCC: data_out = 8'h87;
                    16'hBBCD: data_out = 8'h88;
                    16'hBBCE: data_out = 8'h89;
                    16'hBBCF: data_out = 8'h8A;
                    16'hBBD0: data_out = 8'h8B;
                    16'hBBD1: data_out = 8'h8C;
                    16'hBBD2: data_out = 8'h8D;
                    16'hBBD3: data_out = 8'h8E;
                    16'hBBD4: data_out = 8'h8F;
                    16'hBBD5: data_out = 8'h90;
                    16'hBBD6: data_out = 8'h91;
                    16'hBBD7: data_out = 8'h92;
                    16'hBBD8: data_out = 8'h93;
                    16'hBBD9: data_out = 8'h94;
                    16'hBBDA: data_out = 8'h95;
                    16'hBBDB: data_out = 8'h96;
                    16'hBBDC: data_out = 8'h97;
                    16'hBBDD: data_out = 8'h98;
                    16'hBBDE: data_out = 8'h99;
                    16'hBBDF: data_out = 8'h9A;
                    16'hBBE0: data_out = 8'h9B;
                    16'hBBE1: data_out = 8'h9C;
                    16'hBBE2: data_out = 8'h9D;
                    16'hBBE3: data_out = 8'h9E;
                    16'hBBE4: data_out = 8'h9F;
                    16'hBBE5: data_out = 8'hA0;
                    16'hBBE6: data_out = 8'hA1;
                    16'hBBE7: data_out = 8'hA2;
                    16'hBBE8: data_out = 8'hA3;
                    16'hBBE9: data_out = 8'hA4;
                    16'hBBEA: data_out = 8'hA5;
                    16'hBBEB: data_out = 8'hA6;
                    16'hBBEC: data_out = 8'hA7;
                    16'hBBED: data_out = 8'hA8;
                    16'hBBEE: data_out = 8'hA9;
                    16'hBBEF: data_out = 8'hAA;
                    16'hBBF0: data_out = 8'hAB;
                    16'hBBF1: data_out = 8'hAC;
                    16'hBBF2: data_out = 8'hAD;
                    16'hBBF3: data_out = 8'hAE;
                    16'hBBF4: data_out = 8'hAF;
                    16'hBBF5: data_out = 8'hB0;
                    16'hBBF6: data_out = 8'hB1;
                    16'hBBF7: data_out = 8'hB2;
                    16'hBBF8: data_out = 8'hB3;
                    16'hBBF9: data_out = 8'hB4;
                    16'hBBFA: data_out = 8'hB5;
                    16'hBBFB: data_out = 8'hB6;
                    16'hBBFC: data_out = 8'hB7;
                    16'hBBFD: data_out = 8'hB8;
                    16'hBBFE: data_out = 8'hB9;
                    16'hBBFF: data_out = 8'hBA;
                    16'hBC00: data_out = 8'hBC;
                    16'hBC01: data_out = 8'hBB;
                    16'hBC02: data_out = 8'hBA;
                    16'hBC03: data_out = 8'hB9;
                    16'hBC04: data_out = 8'hB8;
                    16'hBC05: data_out = 8'hB7;
                    16'hBC06: data_out = 8'hB6;
                    16'hBC07: data_out = 8'hB5;
                    16'hBC08: data_out = 8'hB4;
                    16'hBC09: data_out = 8'hB3;
                    16'hBC0A: data_out = 8'hB2;
                    16'hBC0B: data_out = 8'hB1;
                    16'hBC0C: data_out = 8'hB0;
                    16'hBC0D: data_out = 8'hAF;
                    16'hBC0E: data_out = 8'hAE;
                    16'hBC0F: data_out = 8'hAD;
                    16'hBC10: data_out = 8'hAC;
                    16'hBC11: data_out = 8'hAB;
                    16'hBC12: data_out = 8'hAA;
                    16'hBC13: data_out = 8'hA9;
                    16'hBC14: data_out = 8'hA8;
                    16'hBC15: data_out = 8'hA7;
                    16'hBC16: data_out = 8'hA6;
                    16'hBC17: data_out = 8'hA5;
                    16'hBC18: data_out = 8'hA4;
                    16'hBC19: data_out = 8'hA3;
                    16'hBC1A: data_out = 8'hA2;
                    16'hBC1B: data_out = 8'hA1;
                    16'hBC1C: data_out = 8'hA0;
                    16'hBC1D: data_out = 8'h9F;
                    16'hBC1E: data_out = 8'h9E;
                    16'hBC1F: data_out = 8'h9D;
                    16'hBC20: data_out = 8'h9C;
                    16'hBC21: data_out = 8'h9B;
                    16'hBC22: data_out = 8'h9A;
                    16'hBC23: data_out = 8'h99;
                    16'hBC24: data_out = 8'h98;
                    16'hBC25: data_out = 8'h97;
                    16'hBC26: data_out = 8'h96;
                    16'hBC27: data_out = 8'h95;
                    16'hBC28: data_out = 8'h94;
                    16'hBC29: data_out = 8'h93;
                    16'hBC2A: data_out = 8'h92;
                    16'hBC2B: data_out = 8'h91;
                    16'hBC2C: data_out = 8'h90;
                    16'hBC2D: data_out = 8'h8F;
                    16'hBC2E: data_out = 8'h8E;
                    16'hBC2F: data_out = 8'h8D;
                    16'hBC30: data_out = 8'h8C;
                    16'hBC31: data_out = 8'h8B;
                    16'hBC32: data_out = 8'h8A;
                    16'hBC33: data_out = 8'h89;
                    16'hBC34: data_out = 8'h88;
                    16'hBC35: data_out = 8'h87;
                    16'hBC36: data_out = 8'h86;
                    16'hBC37: data_out = 8'h85;
                    16'hBC38: data_out = 8'h84;
                    16'hBC39: data_out = 8'h83;
                    16'hBC3A: data_out = 8'h82;
                    16'hBC3B: data_out = 8'h81;
                    16'hBC3C: data_out = 8'h0;
                    16'hBC3D: data_out = 8'h1;
                    16'hBC3E: data_out = 8'h2;
                    16'hBC3F: data_out = 8'h3;
                    16'hBC40: data_out = 8'h4;
                    16'hBC41: data_out = 8'h5;
                    16'hBC42: data_out = 8'h6;
                    16'hBC43: data_out = 8'h7;
                    16'hBC44: data_out = 8'h8;
                    16'hBC45: data_out = 8'h9;
                    16'hBC46: data_out = 8'hA;
                    16'hBC47: data_out = 8'hB;
                    16'hBC48: data_out = 8'hC;
                    16'hBC49: data_out = 8'hD;
                    16'hBC4A: data_out = 8'hE;
                    16'hBC4B: data_out = 8'hF;
                    16'hBC4C: data_out = 8'h10;
                    16'hBC4D: data_out = 8'h11;
                    16'hBC4E: data_out = 8'h12;
                    16'hBC4F: data_out = 8'h13;
                    16'hBC50: data_out = 8'h14;
                    16'hBC51: data_out = 8'h15;
                    16'hBC52: data_out = 8'h16;
                    16'hBC53: data_out = 8'h17;
                    16'hBC54: data_out = 8'h18;
                    16'hBC55: data_out = 8'h19;
                    16'hBC56: data_out = 8'h1A;
                    16'hBC57: data_out = 8'h1B;
                    16'hBC58: data_out = 8'h1C;
                    16'hBC59: data_out = 8'h1D;
                    16'hBC5A: data_out = 8'h1E;
                    16'hBC5B: data_out = 8'h1F;
                    16'hBC5C: data_out = 8'h20;
                    16'hBC5D: data_out = 8'h21;
                    16'hBC5E: data_out = 8'h22;
                    16'hBC5F: data_out = 8'h23;
                    16'hBC60: data_out = 8'h24;
                    16'hBC61: data_out = 8'h25;
                    16'hBC62: data_out = 8'h26;
                    16'hBC63: data_out = 8'h27;
                    16'hBC64: data_out = 8'h28;
                    16'hBC65: data_out = 8'h29;
                    16'hBC66: data_out = 8'h2A;
                    16'hBC67: data_out = 8'h2B;
                    16'hBC68: data_out = 8'h2C;
                    16'hBC69: data_out = 8'h2D;
                    16'hBC6A: data_out = 8'h2E;
                    16'hBC6B: data_out = 8'h2F;
                    16'hBC6C: data_out = 8'h30;
                    16'hBC6D: data_out = 8'h31;
                    16'hBC6E: data_out = 8'h32;
                    16'hBC6F: data_out = 8'h33;
                    16'hBC70: data_out = 8'h34;
                    16'hBC71: data_out = 8'h35;
                    16'hBC72: data_out = 8'h36;
                    16'hBC73: data_out = 8'h37;
                    16'hBC74: data_out = 8'h38;
                    16'hBC75: data_out = 8'h39;
                    16'hBC76: data_out = 8'h3A;
                    16'hBC77: data_out = 8'h3B;
                    16'hBC78: data_out = 8'h3C;
                    16'hBC79: data_out = 8'h3D;
                    16'hBC7A: data_out = 8'h3E;
                    16'hBC7B: data_out = 8'h3F;
                    16'hBC7C: data_out = 8'h40;
                    16'hBC7D: data_out = 8'h41;
                    16'hBC7E: data_out = 8'h42;
                    16'hBC7F: data_out = 8'h43;
                    16'hBC80: data_out = 8'hBC;
                    16'hBC81: data_out = 8'hBD;
                    16'hBC82: data_out = 8'hBE;
                    16'hBC83: data_out = 8'hBF;
                    16'hBC84: data_out = 8'hC0;
                    16'hBC85: data_out = 8'hC1;
                    16'hBC86: data_out = 8'hC2;
                    16'hBC87: data_out = 8'hC3;
                    16'hBC88: data_out = 8'hC4;
                    16'hBC89: data_out = 8'hC5;
                    16'hBC8A: data_out = 8'hC6;
                    16'hBC8B: data_out = 8'hC7;
                    16'hBC8C: data_out = 8'hC8;
                    16'hBC8D: data_out = 8'hC9;
                    16'hBC8E: data_out = 8'hCA;
                    16'hBC8F: data_out = 8'hCB;
                    16'hBC90: data_out = 8'hCC;
                    16'hBC91: data_out = 8'hCD;
                    16'hBC92: data_out = 8'hCE;
                    16'hBC93: data_out = 8'hCF;
                    16'hBC94: data_out = 8'hD0;
                    16'hBC95: data_out = 8'hD1;
                    16'hBC96: data_out = 8'hD2;
                    16'hBC97: data_out = 8'hD3;
                    16'hBC98: data_out = 8'hD4;
                    16'hBC99: data_out = 8'hD5;
                    16'hBC9A: data_out = 8'hD6;
                    16'hBC9B: data_out = 8'hD7;
                    16'hBC9C: data_out = 8'hD8;
                    16'hBC9D: data_out = 8'hD9;
                    16'hBC9E: data_out = 8'hDA;
                    16'hBC9F: data_out = 8'hDB;
                    16'hBCA0: data_out = 8'hDC;
                    16'hBCA1: data_out = 8'hDD;
                    16'hBCA2: data_out = 8'hDE;
                    16'hBCA3: data_out = 8'hDF;
                    16'hBCA4: data_out = 8'hE0;
                    16'hBCA5: data_out = 8'hE1;
                    16'hBCA6: data_out = 8'hE2;
                    16'hBCA7: data_out = 8'hE3;
                    16'hBCA8: data_out = 8'hE4;
                    16'hBCA9: data_out = 8'hE5;
                    16'hBCAA: data_out = 8'hE6;
                    16'hBCAB: data_out = 8'hE7;
                    16'hBCAC: data_out = 8'hE8;
                    16'hBCAD: data_out = 8'hE9;
                    16'hBCAE: data_out = 8'hEA;
                    16'hBCAF: data_out = 8'hEB;
                    16'hBCB0: data_out = 8'hEC;
                    16'hBCB1: data_out = 8'hED;
                    16'hBCB2: data_out = 8'hEE;
                    16'hBCB3: data_out = 8'hEF;
                    16'hBCB4: data_out = 8'hF0;
                    16'hBCB5: data_out = 8'hF1;
                    16'hBCB6: data_out = 8'hF2;
                    16'hBCB7: data_out = 8'hF3;
                    16'hBCB8: data_out = 8'hF4;
                    16'hBCB9: data_out = 8'hF5;
                    16'hBCBA: data_out = 8'hF6;
                    16'hBCBB: data_out = 8'hF7;
                    16'hBCBC: data_out = 8'hF8;
                    16'hBCBD: data_out = 8'hF9;
                    16'hBCBE: data_out = 8'hFA;
                    16'hBCBF: data_out = 8'hFB;
                    16'hBCC0: data_out = 8'hFC;
                    16'hBCC1: data_out = 8'hFD;
                    16'hBCC2: data_out = 8'hFE;
                    16'hBCC3: data_out = 8'hFF;
                    16'hBCC4: data_out = 8'h80;
                    16'hBCC5: data_out = 8'h81;
                    16'hBCC6: data_out = 8'h82;
                    16'hBCC7: data_out = 8'h83;
                    16'hBCC8: data_out = 8'h84;
                    16'hBCC9: data_out = 8'h85;
                    16'hBCCA: data_out = 8'h86;
                    16'hBCCB: data_out = 8'h87;
                    16'hBCCC: data_out = 8'h88;
                    16'hBCCD: data_out = 8'h89;
                    16'hBCCE: data_out = 8'h8A;
                    16'hBCCF: data_out = 8'h8B;
                    16'hBCD0: data_out = 8'h8C;
                    16'hBCD1: data_out = 8'h8D;
                    16'hBCD2: data_out = 8'h8E;
                    16'hBCD3: data_out = 8'h8F;
                    16'hBCD4: data_out = 8'h90;
                    16'hBCD5: data_out = 8'h91;
                    16'hBCD6: data_out = 8'h92;
                    16'hBCD7: data_out = 8'h93;
                    16'hBCD8: data_out = 8'h94;
                    16'hBCD9: data_out = 8'h95;
                    16'hBCDA: data_out = 8'h96;
                    16'hBCDB: data_out = 8'h97;
                    16'hBCDC: data_out = 8'h98;
                    16'hBCDD: data_out = 8'h99;
                    16'hBCDE: data_out = 8'h9A;
                    16'hBCDF: data_out = 8'h9B;
                    16'hBCE0: data_out = 8'h9C;
                    16'hBCE1: data_out = 8'h9D;
                    16'hBCE2: data_out = 8'h9E;
                    16'hBCE3: data_out = 8'h9F;
                    16'hBCE4: data_out = 8'hA0;
                    16'hBCE5: data_out = 8'hA1;
                    16'hBCE6: data_out = 8'hA2;
                    16'hBCE7: data_out = 8'hA3;
                    16'hBCE8: data_out = 8'hA4;
                    16'hBCE9: data_out = 8'hA5;
                    16'hBCEA: data_out = 8'hA6;
                    16'hBCEB: data_out = 8'hA7;
                    16'hBCEC: data_out = 8'hA8;
                    16'hBCED: data_out = 8'hA9;
                    16'hBCEE: data_out = 8'hAA;
                    16'hBCEF: data_out = 8'hAB;
                    16'hBCF0: data_out = 8'hAC;
                    16'hBCF1: data_out = 8'hAD;
                    16'hBCF2: data_out = 8'hAE;
                    16'hBCF3: data_out = 8'hAF;
                    16'hBCF4: data_out = 8'hB0;
                    16'hBCF5: data_out = 8'hB1;
                    16'hBCF6: data_out = 8'hB2;
                    16'hBCF7: data_out = 8'hB3;
                    16'hBCF8: data_out = 8'hB4;
                    16'hBCF9: data_out = 8'hB5;
                    16'hBCFA: data_out = 8'hB6;
                    16'hBCFB: data_out = 8'hB7;
                    16'hBCFC: data_out = 8'hB8;
                    16'hBCFD: data_out = 8'hB9;
                    16'hBCFE: data_out = 8'hBA;
                    16'hBCFF: data_out = 8'hBB;
                    16'hBD00: data_out = 8'hBD;
                    16'hBD01: data_out = 8'hBC;
                    16'hBD02: data_out = 8'hBB;
                    16'hBD03: data_out = 8'hBA;
                    16'hBD04: data_out = 8'hB9;
                    16'hBD05: data_out = 8'hB8;
                    16'hBD06: data_out = 8'hB7;
                    16'hBD07: data_out = 8'hB6;
                    16'hBD08: data_out = 8'hB5;
                    16'hBD09: data_out = 8'hB4;
                    16'hBD0A: data_out = 8'hB3;
                    16'hBD0B: data_out = 8'hB2;
                    16'hBD0C: data_out = 8'hB1;
                    16'hBD0D: data_out = 8'hB0;
                    16'hBD0E: data_out = 8'hAF;
                    16'hBD0F: data_out = 8'hAE;
                    16'hBD10: data_out = 8'hAD;
                    16'hBD11: data_out = 8'hAC;
                    16'hBD12: data_out = 8'hAB;
                    16'hBD13: data_out = 8'hAA;
                    16'hBD14: data_out = 8'hA9;
                    16'hBD15: data_out = 8'hA8;
                    16'hBD16: data_out = 8'hA7;
                    16'hBD17: data_out = 8'hA6;
                    16'hBD18: data_out = 8'hA5;
                    16'hBD19: data_out = 8'hA4;
                    16'hBD1A: data_out = 8'hA3;
                    16'hBD1B: data_out = 8'hA2;
                    16'hBD1C: data_out = 8'hA1;
                    16'hBD1D: data_out = 8'hA0;
                    16'hBD1E: data_out = 8'h9F;
                    16'hBD1F: data_out = 8'h9E;
                    16'hBD20: data_out = 8'h9D;
                    16'hBD21: data_out = 8'h9C;
                    16'hBD22: data_out = 8'h9B;
                    16'hBD23: data_out = 8'h9A;
                    16'hBD24: data_out = 8'h99;
                    16'hBD25: data_out = 8'h98;
                    16'hBD26: data_out = 8'h97;
                    16'hBD27: data_out = 8'h96;
                    16'hBD28: data_out = 8'h95;
                    16'hBD29: data_out = 8'h94;
                    16'hBD2A: data_out = 8'h93;
                    16'hBD2B: data_out = 8'h92;
                    16'hBD2C: data_out = 8'h91;
                    16'hBD2D: data_out = 8'h90;
                    16'hBD2E: data_out = 8'h8F;
                    16'hBD2F: data_out = 8'h8E;
                    16'hBD30: data_out = 8'h8D;
                    16'hBD31: data_out = 8'h8C;
                    16'hBD32: data_out = 8'h8B;
                    16'hBD33: data_out = 8'h8A;
                    16'hBD34: data_out = 8'h89;
                    16'hBD35: data_out = 8'h88;
                    16'hBD36: data_out = 8'h87;
                    16'hBD37: data_out = 8'h86;
                    16'hBD38: data_out = 8'h85;
                    16'hBD39: data_out = 8'h84;
                    16'hBD3A: data_out = 8'h83;
                    16'hBD3B: data_out = 8'h82;
                    16'hBD3C: data_out = 8'h81;
                    16'hBD3D: data_out = 8'h0;
                    16'hBD3E: data_out = 8'h1;
                    16'hBD3F: data_out = 8'h2;
                    16'hBD40: data_out = 8'h3;
                    16'hBD41: data_out = 8'h4;
                    16'hBD42: data_out = 8'h5;
                    16'hBD43: data_out = 8'h6;
                    16'hBD44: data_out = 8'h7;
                    16'hBD45: data_out = 8'h8;
                    16'hBD46: data_out = 8'h9;
                    16'hBD47: data_out = 8'hA;
                    16'hBD48: data_out = 8'hB;
                    16'hBD49: data_out = 8'hC;
                    16'hBD4A: data_out = 8'hD;
                    16'hBD4B: data_out = 8'hE;
                    16'hBD4C: data_out = 8'hF;
                    16'hBD4D: data_out = 8'h10;
                    16'hBD4E: data_out = 8'h11;
                    16'hBD4F: data_out = 8'h12;
                    16'hBD50: data_out = 8'h13;
                    16'hBD51: data_out = 8'h14;
                    16'hBD52: data_out = 8'h15;
                    16'hBD53: data_out = 8'h16;
                    16'hBD54: data_out = 8'h17;
                    16'hBD55: data_out = 8'h18;
                    16'hBD56: data_out = 8'h19;
                    16'hBD57: data_out = 8'h1A;
                    16'hBD58: data_out = 8'h1B;
                    16'hBD59: data_out = 8'h1C;
                    16'hBD5A: data_out = 8'h1D;
                    16'hBD5B: data_out = 8'h1E;
                    16'hBD5C: data_out = 8'h1F;
                    16'hBD5D: data_out = 8'h20;
                    16'hBD5E: data_out = 8'h21;
                    16'hBD5F: data_out = 8'h22;
                    16'hBD60: data_out = 8'h23;
                    16'hBD61: data_out = 8'h24;
                    16'hBD62: data_out = 8'h25;
                    16'hBD63: data_out = 8'h26;
                    16'hBD64: data_out = 8'h27;
                    16'hBD65: data_out = 8'h28;
                    16'hBD66: data_out = 8'h29;
                    16'hBD67: data_out = 8'h2A;
                    16'hBD68: data_out = 8'h2B;
                    16'hBD69: data_out = 8'h2C;
                    16'hBD6A: data_out = 8'h2D;
                    16'hBD6B: data_out = 8'h2E;
                    16'hBD6C: data_out = 8'h2F;
                    16'hBD6D: data_out = 8'h30;
                    16'hBD6E: data_out = 8'h31;
                    16'hBD6F: data_out = 8'h32;
                    16'hBD70: data_out = 8'h33;
                    16'hBD71: data_out = 8'h34;
                    16'hBD72: data_out = 8'h35;
                    16'hBD73: data_out = 8'h36;
                    16'hBD74: data_out = 8'h37;
                    16'hBD75: data_out = 8'h38;
                    16'hBD76: data_out = 8'h39;
                    16'hBD77: data_out = 8'h3A;
                    16'hBD78: data_out = 8'h3B;
                    16'hBD79: data_out = 8'h3C;
                    16'hBD7A: data_out = 8'h3D;
                    16'hBD7B: data_out = 8'h3E;
                    16'hBD7C: data_out = 8'h3F;
                    16'hBD7D: data_out = 8'h40;
                    16'hBD7E: data_out = 8'h41;
                    16'hBD7F: data_out = 8'h42;
                    16'hBD80: data_out = 8'hBD;
                    16'hBD81: data_out = 8'hBE;
                    16'hBD82: data_out = 8'hBF;
                    16'hBD83: data_out = 8'hC0;
                    16'hBD84: data_out = 8'hC1;
                    16'hBD85: data_out = 8'hC2;
                    16'hBD86: data_out = 8'hC3;
                    16'hBD87: data_out = 8'hC4;
                    16'hBD88: data_out = 8'hC5;
                    16'hBD89: data_out = 8'hC6;
                    16'hBD8A: data_out = 8'hC7;
                    16'hBD8B: data_out = 8'hC8;
                    16'hBD8C: data_out = 8'hC9;
                    16'hBD8D: data_out = 8'hCA;
                    16'hBD8E: data_out = 8'hCB;
                    16'hBD8F: data_out = 8'hCC;
                    16'hBD90: data_out = 8'hCD;
                    16'hBD91: data_out = 8'hCE;
                    16'hBD92: data_out = 8'hCF;
                    16'hBD93: data_out = 8'hD0;
                    16'hBD94: data_out = 8'hD1;
                    16'hBD95: data_out = 8'hD2;
                    16'hBD96: data_out = 8'hD3;
                    16'hBD97: data_out = 8'hD4;
                    16'hBD98: data_out = 8'hD5;
                    16'hBD99: data_out = 8'hD6;
                    16'hBD9A: data_out = 8'hD7;
                    16'hBD9B: data_out = 8'hD8;
                    16'hBD9C: data_out = 8'hD9;
                    16'hBD9D: data_out = 8'hDA;
                    16'hBD9E: data_out = 8'hDB;
                    16'hBD9F: data_out = 8'hDC;
                    16'hBDA0: data_out = 8'hDD;
                    16'hBDA1: data_out = 8'hDE;
                    16'hBDA2: data_out = 8'hDF;
                    16'hBDA3: data_out = 8'hE0;
                    16'hBDA4: data_out = 8'hE1;
                    16'hBDA5: data_out = 8'hE2;
                    16'hBDA6: data_out = 8'hE3;
                    16'hBDA7: data_out = 8'hE4;
                    16'hBDA8: data_out = 8'hE5;
                    16'hBDA9: data_out = 8'hE6;
                    16'hBDAA: data_out = 8'hE7;
                    16'hBDAB: data_out = 8'hE8;
                    16'hBDAC: data_out = 8'hE9;
                    16'hBDAD: data_out = 8'hEA;
                    16'hBDAE: data_out = 8'hEB;
                    16'hBDAF: data_out = 8'hEC;
                    16'hBDB0: data_out = 8'hED;
                    16'hBDB1: data_out = 8'hEE;
                    16'hBDB2: data_out = 8'hEF;
                    16'hBDB3: data_out = 8'hF0;
                    16'hBDB4: data_out = 8'hF1;
                    16'hBDB5: data_out = 8'hF2;
                    16'hBDB6: data_out = 8'hF3;
                    16'hBDB7: data_out = 8'hF4;
                    16'hBDB8: data_out = 8'hF5;
                    16'hBDB9: data_out = 8'hF6;
                    16'hBDBA: data_out = 8'hF7;
                    16'hBDBB: data_out = 8'hF8;
                    16'hBDBC: data_out = 8'hF9;
                    16'hBDBD: data_out = 8'hFA;
                    16'hBDBE: data_out = 8'hFB;
                    16'hBDBF: data_out = 8'hFC;
                    16'hBDC0: data_out = 8'hFD;
                    16'hBDC1: data_out = 8'hFE;
                    16'hBDC2: data_out = 8'hFF;
                    16'hBDC3: data_out = 8'h80;
                    16'hBDC4: data_out = 8'h81;
                    16'hBDC5: data_out = 8'h82;
                    16'hBDC6: data_out = 8'h83;
                    16'hBDC7: data_out = 8'h84;
                    16'hBDC8: data_out = 8'h85;
                    16'hBDC9: data_out = 8'h86;
                    16'hBDCA: data_out = 8'h87;
                    16'hBDCB: data_out = 8'h88;
                    16'hBDCC: data_out = 8'h89;
                    16'hBDCD: data_out = 8'h8A;
                    16'hBDCE: data_out = 8'h8B;
                    16'hBDCF: data_out = 8'h8C;
                    16'hBDD0: data_out = 8'h8D;
                    16'hBDD1: data_out = 8'h8E;
                    16'hBDD2: data_out = 8'h8F;
                    16'hBDD3: data_out = 8'h90;
                    16'hBDD4: data_out = 8'h91;
                    16'hBDD5: data_out = 8'h92;
                    16'hBDD6: data_out = 8'h93;
                    16'hBDD7: data_out = 8'h94;
                    16'hBDD8: data_out = 8'h95;
                    16'hBDD9: data_out = 8'h96;
                    16'hBDDA: data_out = 8'h97;
                    16'hBDDB: data_out = 8'h98;
                    16'hBDDC: data_out = 8'h99;
                    16'hBDDD: data_out = 8'h9A;
                    16'hBDDE: data_out = 8'h9B;
                    16'hBDDF: data_out = 8'h9C;
                    16'hBDE0: data_out = 8'h9D;
                    16'hBDE1: data_out = 8'h9E;
                    16'hBDE2: data_out = 8'h9F;
                    16'hBDE3: data_out = 8'hA0;
                    16'hBDE4: data_out = 8'hA1;
                    16'hBDE5: data_out = 8'hA2;
                    16'hBDE6: data_out = 8'hA3;
                    16'hBDE7: data_out = 8'hA4;
                    16'hBDE8: data_out = 8'hA5;
                    16'hBDE9: data_out = 8'hA6;
                    16'hBDEA: data_out = 8'hA7;
                    16'hBDEB: data_out = 8'hA8;
                    16'hBDEC: data_out = 8'hA9;
                    16'hBDED: data_out = 8'hAA;
                    16'hBDEE: data_out = 8'hAB;
                    16'hBDEF: data_out = 8'hAC;
                    16'hBDF0: data_out = 8'hAD;
                    16'hBDF1: data_out = 8'hAE;
                    16'hBDF2: data_out = 8'hAF;
                    16'hBDF3: data_out = 8'hB0;
                    16'hBDF4: data_out = 8'hB1;
                    16'hBDF5: data_out = 8'hB2;
                    16'hBDF6: data_out = 8'hB3;
                    16'hBDF7: data_out = 8'hB4;
                    16'hBDF8: data_out = 8'hB5;
                    16'hBDF9: data_out = 8'hB6;
                    16'hBDFA: data_out = 8'hB7;
                    16'hBDFB: data_out = 8'hB8;
                    16'hBDFC: data_out = 8'hB9;
                    16'hBDFD: data_out = 8'hBA;
                    16'hBDFE: data_out = 8'hBB;
                    16'hBDFF: data_out = 8'hBC;
                    16'hBE00: data_out = 8'hBE;
                    16'hBE01: data_out = 8'hBD;
                    16'hBE02: data_out = 8'hBC;
                    16'hBE03: data_out = 8'hBB;
                    16'hBE04: data_out = 8'hBA;
                    16'hBE05: data_out = 8'hB9;
                    16'hBE06: data_out = 8'hB8;
                    16'hBE07: data_out = 8'hB7;
                    16'hBE08: data_out = 8'hB6;
                    16'hBE09: data_out = 8'hB5;
                    16'hBE0A: data_out = 8'hB4;
                    16'hBE0B: data_out = 8'hB3;
                    16'hBE0C: data_out = 8'hB2;
                    16'hBE0D: data_out = 8'hB1;
                    16'hBE0E: data_out = 8'hB0;
                    16'hBE0F: data_out = 8'hAF;
                    16'hBE10: data_out = 8'hAE;
                    16'hBE11: data_out = 8'hAD;
                    16'hBE12: data_out = 8'hAC;
                    16'hBE13: data_out = 8'hAB;
                    16'hBE14: data_out = 8'hAA;
                    16'hBE15: data_out = 8'hA9;
                    16'hBE16: data_out = 8'hA8;
                    16'hBE17: data_out = 8'hA7;
                    16'hBE18: data_out = 8'hA6;
                    16'hBE19: data_out = 8'hA5;
                    16'hBE1A: data_out = 8'hA4;
                    16'hBE1B: data_out = 8'hA3;
                    16'hBE1C: data_out = 8'hA2;
                    16'hBE1D: data_out = 8'hA1;
                    16'hBE1E: data_out = 8'hA0;
                    16'hBE1F: data_out = 8'h9F;
                    16'hBE20: data_out = 8'h9E;
                    16'hBE21: data_out = 8'h9D;
                    16'hBE22: data_out = 8'h9C;
                    16'hBE23: data_out = 8'h9B;
                    16'hBE24: data_out = 8'h9A;
                    16'hBE25: data_out = 8'h99;
                    16'hBE26: data_out = 8'h98;
                    16'hBE27: data_out = 8'h97;
                    16'hBE28: data_out = 8'h96;
                    16'hBE29: data_out = 8'h95;
                    16'hBE2A: data_out = 8'h94;
                    16'hBE2B: data_out = 8'h93;
                    16'hBE2C: data_out = 8'h92;
                    16'hBE2D: data_out = 8'h91;
                    16'hBE2E: data_out = 8'h90;
                    16'hBE2F: data_out = 8'h8F;
                    16'hBE30: data_out = 8'h8E;
                    16'hBE31: data_out = 8'h8D;
                    16'hBE32: data_out = 8'h8C;
                    16'hBE33: data_out = 8'h8B;
                    16'hBE34: data_out = 8'h8A;
                    16'hBE35: data_out = 8'h89;
                    16'hBE36: data_out = 8'h88;
                    16'hBE37: data_out = 8'h87;
                    16'hBE38: data_out = 8'h86;
                    16'hBE39: data_out = 8'h85;
                    16'hBE3A: data_out = 8'h84;
                    16'hBE3B: data_out = 8'h83;
                    16'hBE3C: data_out = 8'h82;
                    16'hBE3D: data_out = 8'h81;
                    16'hBE3E: data_out = 8'h0;
                    16'hBE3F: data_out = 8'h1;
                    16'hBE40: data_out = 8'h2;
                    16'hBE41: data_out = 8'h3;
                    16'hBE42: data_out = 8'h4;
                    16'hBE43: data_out = 8'h5;
                    16'hBE44: data_out = 8'h6;
                    16'hBE45: data_out = 8'h7;
                    16'hBE46: data_out = 8'h8;
                    16'hBE47: data_out = 8'h9;
                    16'hBE48: data_out = 8'hA;
                    16'hBE49: data_out = 8'hB;
                    16'hBE4A: data_out = 8'hC;
                    16'hBE4B: data_out = 8'hD;
                    16'hBE4C: data_out = 8'hE;
                    16'hBE4D: data_out = 8'hF;
                    16'hBE4E: data_out = 8'h10;
                    16'hBE4F: data_out = 8'h11;
                    16'hBE50: data_out = 8'h12;
                    16'hBE51: data_out = 8'h13;
                    16'hBE52: data_out = 8'h14;
                    16'hBE53: data_out = 8'h15;
                    16'hBE54: data_out = 8'h16;
                    16'hBE55: data_out = 8'h17;
                    16'hBE56: data_out = 8'h18;
                    16'hBE57: data_out = 8'h19;
                    16'hBE58: data_out = 8'h1A;
                    16'hBE59: data_out = 8'h1B;
                    16'hBE5A: data_out = 8'h1C;
                    16'hBE5B: data_out = 8'h1D;
                    16'hBE5C: data_out = 8'h1E;
                    16'hBE5D: data_out = 8'h1F;
                    16'hBE5E: data_out = 8'h20;
                    16'hBE5F: data_out = 8'h21;
                    16'hBE60: data_out = 8'h22;
                    16'hBE61: data_out = 8'h23;
                    16'hBE62: data_out = 8'h24;
                    16'hBE63: data_out = 8'h25;
                    16'hBE64: data_out = 8'h26;
                    16'hBE65: data_out = 8'h27;
                    16'hBE66: data_out = 8'h28;
                    16'hBE67: data_out = 8'h29;
                    16'hBE68: data_out = 8'h2A;
                    16'hBE69: data_out = 8'h2B;
                    16'hBE6A: data_out = 8'h2C;
                    16'hBE6B: data_out = 8'h2D;
                    16'hBE6C: data_out = 8'h2E;
                    16'hBE6D: data_out = 8'h2F;
                    16'hBE6E: data_out = 8'h30;
                    16'hBE6F: data_out = 8'h31;
                    16'hBE70: data_out = 8'h32;
                    16'hBE71: data_out = 8'h33;
                    16'hBE72: data_out = 8'h34;
                    16'hBE73: data_out = 8'h35;
                    16'hBE74: data_out = 8'h36;
                    16'hBE75: data_out = 8'h37;
                    16'hBE76: data_out = 8'h38;
                    16'hBE77: data_out = 8'h39;
                    16'hBE78: data_out = 8'h3A;
                    16'hBE79: data_out = 8'h3B;
                    16'hBE7A: data_out = 8'h3C;
                    16'hBE7B: data_out = 8'h3D;
                    16'hBE7C: data_out = 8'h3E;
                    16'hBE7D: data_out = 8'h3F;
                    16'hBE7E: data_out = 8'h40;
                    16'hBE7F: data_out = 8'h41;
                    16'hBE80: data_out = 8'hBE;
                    16'hBE81: data_out = 8'hBF;
                    16'hBE82: data_out = 8'hC0;
                    16'hBE83: data_out = 8'hC1;
                    16'hBE84: data_out = 8'hC2;
                    16'hBE85: data_out = 8'hC3;
                    16'hBE86: data_out = 8'hC4;
                    16'hBE87: data_out = 8'hC5;
                    16'hBE88: data_out = 8'hC6;
                    16'hBE89: data_out = 8'hC7;
                    16'hBE8A: data_out = 8'hC8;
                    16'hBE8B: data_out = 8'hC9;
                    16'hBE8C: data_out = 8'hCA;
                    16'hBE8D: data_out = 8'hCB;
                    16'hBE8E: data_out = 8'hCC;
                    16'hBE8F: data_out = 8'hCD;
                    16'hBE90: data_out = 8'hCE;
                    16'hBE91: data_out = 8'hCF;
                    16'hBE92: data_out = 8'hD0;
                    16'hBE93: data_out = 8'hD1;
                    16'hBE94: data_out = 8'hD2;
                    16'hBE95: data_out = 8'hD3;
                    16'hBE96: data_out = 8'hD4;
                    16'hBE97: data_out = 8'hD5;
                    16'hBE98: data_out = 8'hD6;
                    16'hBE99: data_out = 8'hD7;
                    16'hBE9A: data_out = 8'hD8;
                    16'hBE9B: data_out = 8'hD9;
                    16'hBE9C: data_out = 8'hDA;
                    16'hBE9D: data_out = 8'hDB;
                    16'hBE9E: data_out = 8'hDC;
                    16'hBE9F: data_out = 8'hDD;
                    16'hBEA0: data_out = 8'hDE;
                    16'hBEA1: data_out = 8'hDF;
                    16'hBEA2: data_out = 8'hE0;
                    16'hBEA3: data_out = 8'hE1;
                    16'hBEA4: data_out = 8'hE2;
                    16'hBEA5: data_out = 8'hE3;
                    16'hBEA6: data_out = 8'hE4;
                    16'hBEA7: data_out = 8'hE5;
                    16'hBEA8: data_out = 8'hE6;
                    16'hBEA9: data_out = 8'hE7;
                    16'hBEAA: data_out = 8'hE8;
                    16'hBEAB: data_out = 8'hE9;
                    16'hBEAC: data_out = 8'hEA;
                    16'hBEAD: data_out = 8'hEB;
                    16'hBEAE: data_out = 8'hEC;
                    16'hBEAF: data_out = 8'hED;
                    16'hBEB0: data_out = 8'hEE;
                    16'hBEB1: data_out = 8'hEF;
                    16'hBEB2: data_out = 8'hF0;
                    16'hBEB3: data_out = 8'hF1;
                    16'hBEB4: data_out = 8'hF2;
                    16'hBEB5: data_out = 8'hF3;
                    16'hBEB6: data_out = 8'hF4;
                    16'hBEB7: data_out = 8'hF5;
                    16'hBEB8: data_out = 8'hF6;
                    16'hBEB9: data_out = 8'hF7;
                    16'hBEBA: data_out = 8'hF8;
                    16'hBEBB: data_out = 8'hF9;
                    16'hBEBC: data_out = 8'hFA;
                    16'hBEBD: data_out = 8'hFB;
                    16'hBEBE: data_out = 8'hFC;
                    16'hBEBF: data_out = 8'hFD;
                    16'hBEC0: data_out = 8'hFE;
                    16'hBEC1: data_out = 8'hFF;
                    16'hBEC2: data_out = 8'h80;
                    16'hBEC3: data_out = 8'h81;
                    16'hBEC4: data_out = 8'h82;
                    16'hBEC5: data_out = 8'h83;
                    16'hBEC6: data_out = 8'h84;
                    16'hBEC7: data_out = 8'h85;
                    16'hBEC8: data_out = 8'h86;
                    16'hBEC9: data_out = 8'h87;
                    16'hBECA: data_out = 8'h88;
                    16'hBECB: data_out = 8'h89;
                    16'hBECC: data_out = 8'h8A;
                    16'hBECD: data_out = 8'h8B;
                    16'hBECE: data_out = 8'h8C;
                    16'hBECF: data_out = 8'h8D;
                    16'hBED0: data_out = 8'h8E;
                    16'hBED1: data_out = 8'h8F;
                    16'hBED2: data_out = 8'h90;
                    16'hBED3: data_out = 8'h91;
                    16'hBED4: data_out = 8'h92;
                    16'hBED5: data_out = 8'h93;
                    16'hBED6: data_out = 8'h94;
                    16'hBED7: data_out = 8'h95;
                    16'hBED8: data_out = 8'h96;
                    16'hBED9: data_out = 8'h97;
                    16'hBEDA: data_out = 8'h98;
                    16'hBEDB: data_out = 8'h99;
                    16'hBEDC: data_out = 8'h9A;
                    16'hBEDD: data_out = 8'h9B;
                    16'hBEDE: data_out = 8'h9C;
                    16'hBEDF: data_out = 8'h9D;
                    16'hBEE0: data_out = 8'h9E;
                    16'hBEE1: data_out = 8'h9F;
                    16'hBEE2: data_out = 8'hA0;
                    16'hBEE3: data_out = 8'hA1;
                    16'hBEE4: data_out = 8'hA2;
                    16'hBEE5: data_out = 8'hA3;
                    16'hBEE6: data_out = 8'hA4;
                    16'hBEE7: data_out = 8'hA5;
                    16'hBEE8: data_out = 8'hA6;
                    16'hBEE9: data_out = 8'hA7;
                    16'hBEEA: data_out = 8'hA8;
                    16'hBEEB: data_out = 8'hA9;
                    16'hBEEC: data_out = 8'hAA;
                    16'hBEED: data_out = 8'hAB;
                    16'hBEEE: data_out = 8'hAC;
                    16'hBEEF: data_out = 8'hAD;
                    16'hBEF0: data_out = 8'hAE;
                    16'hBEF1: data_out = 8'hAF;
                    16'hBEF2: data_out = 8'hB0;
                    16'hBEF3: data_out = 8'hB1;
                    16'hBEF4: data_out = 8'hB2;
                    16'hBEF5: data_out = 8'hB3;
                    16'hBEF6: data_out = 8'hB4;
                    16'hBEF7: data_out = 8'hB5;
                    16'hBEF8: data_out = 8'hB6;
                    16'hBEF9: data_out = 8'hB7;
                    16'hBEFA: data_out = 8'hB8;
                    16'hBEFB: data_out = 8'hB9;
                    16'hBEFC: data_out = 8'hBA;
                    16'hBEFD: data_out = 8'hBB;
                    16'hBEFE: data_out = 8'hBC;
                    16'hBEFF: data_out = 8'hBD;
                    16'hBF00: data_out = 8'hBF;
                    16'hBF01: data_out = 8'hBE;
                    16'hBF02: data_out = 8'hBD;
                    16'hBF03: data_out = 8'hBC;
                    16'hBF04: data_out = 8'hBB;
                    16'hBF05: data_out = 8'hBA;
                    16'hBF06: data_out = 8'hB9;
                    16'hBF07: data_out = 8'hB8;
                    16'hBF08: data_out = 8'hB7;
                    16'hBF09: data_out = 8'hB6;
                    16'hBF0A: data_out = 8'hB5;
                    16'hBF0B: data_out = 8'hB4;
                    16'hBF0C: data_out = 8'hB3;
                    16'hBF0D: data_out = 8'hB2;
                    16'hBF0E: data_out = 8'hB1;
                    16'hBF0F: data_out = 8'hB0;
                    16'hBF10: data_out = 8'hAF;
                    16'hBF11: data_out = 8'hAE;
                    16'hBF12: data_out = 8'hAD;
                    16'hBF13: data_out = 8'hAC;
                    16'hBF14: data_out = 8'hAB;
                    16'hBF15: data_out = 8'hAA;
                    16'hBF16: data_out = 8'hA9;
                    16'hBF17: data_out = 8'hA8;
                    16'hBF18: data_out = 8'hA7;
                    16'hBF19: data_out = 8'hA6;
                    16'hBF1A: data_out = 8'hA5;
                    16'hBF1B: data_out = 8'hA4;
                    16'hBF1C: data_out = 8'hA3;
                    16'hBF1D: data_out = 8'hA2;
                    16'hBF1E: data_out = 8'hA1;
                    16'hBF1F: data_out = 8'hA0;
                    16'hBF20: data_out = 8'h9F;
                    16'hBF21: data_out = 8'h9E;
                    16'hBF22: data_out = 8'h9D;
                    16'hBF23: data_out = 8'h9C;
                    16'hBF24: data_out = 8'h9B;
                    16'hBF25: data_out = 8'h9A;
                    16'hBF26: data_out = 8'h99;
                    16'hBF27: data_out = 8'h98;
                    16'hBF28: data_out = 8'h97;
                    16'hBF29: data_out = 8'h96;
                    16'hBF2A: data_out = 8'h95;
                    16'hBF2B: data_out = 8'h94;
                    16'hBF2C: data_out = 8'h93;
                    16'hBF2D: data_out = 8'h92;
                    16'hBF2E: data_out = 8'h91;
                    16'hBF2F: data_out = 8'h90;
                    16'hBF30: data_out = 8'h8F;
                    16'hBF31: data_out = 8'h8E;
                    16'hBF32: data_out = 8'h8D;
                    16'hBF33: data_out = 8'h8C;
                    16'hBF34: data_out = 8'h8B;
                    16'hBF35: data_out = 8'h8A;
                    16'hBF36: data_out = 8'h89;
                    16'hBF37: data_out = 8'h88;
                    16'hBF38: data_out = 8'h87;
                    16'hBF39: data_out = 8'h86;
                    16'hBF3A: data_out = 8'h85;
                    16'hBF3B: data_out = 8'h84;
                    16'hBF3C: data_out = 8'h83;
                    16'hBF3D: data_out = 8'h82;
                    16'hBF3E: data_out = 8'h81;
                    16'hBF3F: data_out = 8'h0;
                    16'hBF40: data_out = 8'h1;
                    16'hBF41: data_out = 8'h2;
                    16'hBF42: data_out = 8'h3;
                    16'hBF43: data_out = 8'h4;
                    16'hBF44: data_out = 8'h5;
                    16'hBF45: data_out = 8'h6;
                    16'hBF46: data_out = 8'h7;
                    16'hBF47: data_out = 8'h8;
                    16'hBF48: data_out = 8'h9;
                    16'hBF49: data_out = 8'hA;
                    16'hBF4A: data_out = 8'hB;
                    16'hBF4B: data_out = 8'hC;
                    16'hBF4C: data_out = 8'hD;
                    16'hBF4D: data_out = 8'hE;
                    16'hBF4E: data_out = 8'hF;
                    16'hBF4F: data_out = 8'h10;
                    16'hBF50: data_out = 8'h11;
                    16'hBF51: data_out = 8'h12;
                    16'hBF52: data_out = 8'h13;
                    16'hBF53: data_out = 8'h14;
                    16'hBF54: data_out = 8'h15;
                    16'hBF55: data_out = 8'h16;
                    16'hBF56: data_out = 8'h17;
                    16'hBF57: data_out = 8'h18;
                    16'hBF58: data_out = 8'h19;
                    16'hBF59: data_out = 8'h1A;
                    16'hBF5A: data_out = 8'h1B;
                    16'hBF5B: data_out = 8'h1C;
                    16'hBF5C: data_out = 8'h1D;
                    16'hBF5D: data_out = 8'h1E;
                    16'hBF5E: data_out = 8'h1F;
                    16'hBF5F: data_out = 8'h20;
                    16'hBF60: data_out = 8'h21;
                    16'hBF61: data_out = 8'h22;
                    16'hBF62: data_out = 8'h23;
                    16'hBF63: data_out = 8'h24;
                    16'hBF64: data_out = 8'h25;
                    16'hBF65: data_out = 8'h26;
                    16'hBF66: data_out = 8'h27;
                    16'hBF67: data_out = 8'h28;
                    16'hBF68: data_out = 8'h29;
                    16'hBF69: data_out = 8'h2A;
                    16'hBF6A: data_out = 8'h2B;
                    16'hBF6B: data_out = 8'h2C;
                    16'hBF6C: data_out = 8'h2D;
                    16'hBF6D: data_out = 8'h2E;
                    16'hBF6E: data_out = 8'h2F;
                    16'hBF6F: data_out = 8'h30;
                    16'hBF70: data_out = 8'h31;
                    16'hBF71: data_out = 8'h32;
                    16'hBF72: data_out = 8'h33;
                    16'hBF73: data_out = 8'h34;
                    16'hBF74: data_out = 8'h35;
                    16'hBF75: data_out = 8'h36;
                    16'hBF76: data_out = 8'h37;
                    16'hBF77: data_out = 8'h38;
                    16'hBF78: data_out = 8'h39;
                    16'hBF79: data_out = 8'h3A;
                    16'hBF7A: data_out = 8'h3B;
                    16'hBF7B: data_out = 8'h3C;
                    16'hBF7C: data_out = 8'h3D;
                    16'hBF7D: data_out = 8'h3E;
                    16'hBF7E: data_out = 8'h3F;
                    16'hBF7F: data_out = 8'h40;
                    16'hBF80: data_out = 8'hBF;
                    16'hBF81: data_out = 8'hC0;
                    16'hBF82: data_out = 8'hC1;
                    16'hBF83: data_out = 8'hC2;
                    16'hBF84: data_out = 8'hC3;
                    16'hBF85: data_out = 8'hC4;
                    16'hBF86: data_out = 8'hC5;
                    16'hBF87: data_out = 8'hC6;
                    16'hBF88: data_out = 8'hC7;
                    16'hBF89: data_out = 8'hC8;
                    16'hBF8A: data_out = 8'hC9;
                    16'hBF8B: data_out = 8'hCA;
                    16'hBF8C: data_out = 8'hCB;
                    16'hBF8D: data_out = 8'hCC;
                    16'hBF8E: data_out = 8'hCD;
                    16'hBF8F: data_out = 8'hCE;
                    16'hBF90: data_out = 8'hCF;
                    16'hBF91: data_out = 8'hD0;
                    16'hBF92: data_out = 8'hD1;
                    16'hBF93: data_out = 8'hD2;
                    16'hBF94: data_out = 8'hD3;
                    16'hBF95: data_out = 8'hD4;
                    16'hBF96: data_out = 8'hD5;
                    16'hBF97: data_out = 8'hD6;
                    16'hBF98: data_out = 8'hD7;
                    16'hBF99: data_out = 8'hD8;
                    16'hBF9A: data_out = 8'hD9;
                    16'hBF9B: data_out = 8'hDA;
                    16'hBF9C: data_out = 8'hDB;
                    16'hBF9D: data_out = 8'hDC;
                    16'hBF9E: data_out = 8'hDD;
                    16'hBF9F: data_out = 8'hDE;
                    16'hBFA0: data_out = 8'hDF;
                    16'hBFA1: data_out = 8'hE0;
                    16'hBFA2: data_out = 8'hE1;
                    16'hBFA3: data_out = 8'hE2;
                    16'hBFA4: data_out = 8'hE3;
                    16'hBFA5: data_out = 8'hE4;
                    16'hBFA6: data_out = 8'hE5;
                    16'hBFA7: data_out = 8'hE6;
                    16'hBFA8: data_out = 8'hE7;
                    16'hBFA9: data_out = 8'hE8;
                    16'hBFAA: data_out = 8'hE9;
                    16'hBFAB: data_out = 8'hEA;
                    16'hBFAC: data_out = 8'hEB;
                    16'hBFAD: data_out = 8'hEC;
                    16'hBFAE: data_out = 8'hED;
                    16'hBFAF: data_out = 8'hEE;
                    16'hBFB0: data_out = 8'hEF;
                    16'hBFB1: data_out = 8'hF0;
                    16'hBFB2: data_out = 8'hF1;
                    16'hBFB3: data_out = 8'hF2;
                    16'hBFB4: data_out = 8'hF3;
                    16'hBFB5: data_out = 8'hF4;
                    16'hBFB6: data_out = 8'hF5;
                    16'hBFB7: data_out = 8'hF6;
                    16'hBFB8: data_out = 8'hF7;
                    16'hBFB9: data_out = 8'hF8;
                    16'hBFBA: data_out = 8'hF9;
                    16'hBFBB: data_out = 8'hFA;
                    16'hBFBC: data_out = 8'hFB;
                    16'hBFBD: data_out = 8'hFC;
                    16'hBFBE: data_out = 8'hFD;
                    16'hBFBF: data_out = 8'hFE;
                    16'hBFC0: data_out = 8'hFF;
                    16'hBFC1: data_out = 8'h80;
                    16'hBFC2: data_out = 8'h81;
                    16'hBFC3: data_out = 8'h82;
                    16'hBFC4: data_out = 8'h83;
                    16'hBFC5: data_out = 8'h84;
                    16'hBFC6: data_out = 8'h85;
                    16'hBFC7: data_out = 8'h86;
                    16'hBFC8: data_out = 8'h87;
                    16'hBFC9: data_out = 8'h88;
                    16'hBFCA: data_out = 8'h89;
                    16'hBFCB: data_out = 8'h8A;
                    16'hBFCC: data_out = 8'h8B;
                    16'hBFCD: data_out = 8'h8C;
                    16'hBFCE: data_out = 8'h8D;
                    16'hBFCF: data_out = 8'h8E;
                    16'hBFD0: data_out = 8'h8F;
                    16'hBFD1: data_out = 8'h90;
                    16'hBFD2: data_out = 8'h91;
                    16'hBFD3: data_out = 8'h92;
                    16'hBFD4: data_out = 8'h93;
                    16'hBFD5: data_out = 8'h94;
                    16'hBFD6: data_out = 8'h95;
                    16'hBFD7: data_out = 8'h96;
                    16'hBFD8: data_out = 8'h97;
                    16'hBFD9: data_out = 8'h98;
                    16'hBFDA: data_out = 8'h99;
                    16'hBFDB: data_out = 8'h9A;
                    16'hBFDC: data_out = 8'h9B;
                    16'hBFDD: data_out = 8'h9C;
                    16'hBFDE: data_out = 8'h9D;
                    16'hBFDF: data_out = 8'h9E;
                    16'hBFE0: data_out = 8'h9F;
                    16'hBFE1: data_out = 8'hA0;
                    16'hBFE2: data_out = 8'hA1;
                    16'hBFE3: data_out = 8'hA2;
                    16'hBFE4: data_out = 8'hA3;
                    16'hBFE5: data_out = 8'hA4;
                    16'hBFE6: data_out = 8'hA5;
                    16'hBFE7: data_out = 8'hA6;
                    16'hBFE8: data_out = 8'hA7;
                    16'hBFE9: data_out = 8'hA8;
                    16'hBFEA: data_out = 8'hA9;
                    16'hBFEB: data_out = 8'hAA;
                    16'hBFEC: data_out = 8'hAB;
                    16'hBFED: data_out = 8'hAC;
                    16'hBFEE: data_out = 8'hAD;
                    16'hBFEF: data_out = 8'hAE;
                    16'hBFF0: data_out = 8'hAF;
                    16'hBFF1: data_out = 8'hB0;
                    16'hBFF2: data_out = 8'hB1;
                    16'hBFF3: data_out = 8'hB2;
                    16'hBFF4: data_out = 8'hB3;
                    16'hBFF5: data_out = 8'hB4;
                    16'hBFF6: data_out = 8'hB5;
                    16'hBFF7: data_out = 8'hB6;
                    16'hBFF8: data_out = 8'hB7;
                    16'hBFF9: data_out = 8'hB8;
                    16'hBFFA: data_out = 8'hB9;
                    16'hBFFB: data_out = 8'hBA;
                    16'hBFFC: data_out = 8'hBB;
                    16'hBFFD: data_out = 8'hBC;
                    16'hBFFE: data_out = 8'hBD;
                    16'hBFFF: data_out = 8'hBE;
                    16'hC000: data_out = 8'hC0;
                    16'hC001: data_out = 8'hBF;
                    16'hC002: data_out = 8'hBE;
                    16'hC003: data_out = 8'hBD;
                    16'hC004: data_out = 8'hBC;
                    16'hC005: data_out = 8'hBB;
                    16'hC006: data_out = 8'hBA;
                    16'hC007: data_out = 8'hB9;
                    16'hC008: data_out = 8'hB8;
                    16'hC009: data_out = 8'hB7;
                    16'hC00A: data_out = 8'hB6;
                    16'hC00B: data_out = 8'hB5;
                    16'hC00C: data_out = 8'hB4;
                    16'hC00D: data_out = 8'hB3;
                    16'hC00E: data_out = 8'hB2;
                    16'hC00F: data_out = 8'hB1;
                    16'hC010: data_out = 8'hB0;
                    16'hC011: data_out = 8'hAF;
                    16'hC012: data_out = 8'hAE;
                    16'hC013: data_out = 8'hAD;
                    16'hC014: data_out = 8'hAC;
                    16'hC015: data_out = 8'hAB;
                    16'hC016: data_out = 8'hAA;
                    16'hC017: data_out = 8'hA9;
                    16'hC018: data_out = 8'hA8;
                    16'hC019: data_out = 8'hA7;
                    16'hC01A: data_out = 8'hA6;
                    16'hC01B: data_out = 8'hA5;
                    16'hC01C: data_out = 8'hA4;
                    16'hC01D: data_out = 8'hA3;
                    16'hC01E: data_out = 8'hA2;
                    16'hC01F: data_out = 8'hA1;
                    16'hC020: data_out = 8'hA0;
                    16'hC021: data_out = 8'h9F;
                    16'hC022: data_out = 8'h9E;
                    16'hC023: data_out = 8'h9D;
                    16'hC024: data_out = 8'h9C;
                    16'hC025: data_out = 8'h9B;
                    16'hC026: data_out = 8'h9A;
                    16'hC027: data_out = 8'h99;
                    16'hC028: data_out = 8'h98;
                    16'hC029: data_out = 8'h97;
                    16'hC02A: data_out = 8'h96;
                    16'hC02B: data_out = 8'h95;
                    16'hC02C: data_out = 8'h94;
                    16'hC02D: data_out = 8'h93;
                    16'hC02E: data_out = 8'h92;
                    16'hC02F: data_out = 8'h91;
                    16'hC030: data_out = 8'h90;
                    16'hC031: data_out = 8'h8F;
                    16'hC032: data_out = 8'h8E;
                    16'hC033: data_out = 8'h8D;
                    16'hC034: data_out = 8'h8C;
                    16'hC035: data_out = 8'h8B;
                    16'hC036: data_out = 8'h8A;
                    16'hC037: data_out = 8'h89;
                    16'hC038: data_out = 8'h88;
                    16'hC039: data_out = 8'h87;
                    16'hC03A: data_out = 8'h86;
                    16'hC03B: data_out = 8'h85;
                    16'hC03C: data_out = 8'h84;
                    16'hC03D: data_out = 8'h83;
                    16'hC03E: data_out = 8'h82;
                    16'hC03F: data_out = 8'h81;
                    16'hC040: data_out = 8'h0;
                    16'hC041: data_out = 8'h1;
                    16'hC042: data_out = 8'h2;
                    16'hC043: data_out = 8'h3;
                    16'hC044: data_out = 8'h4;
                    16'hC045: data_out = 8'h5;
                    16'hC046: data_out = 8'h6;
                    16'hC047: data_out = 8'h7;
                    16'hC048: data_out = 8'h8;
                    16'hC049: data_out = 8'h9;
                    16'hC04A: data_out = 8'hA;
                    16'hC04B: data_out = 8'hB;
                    16'hC04C: data_out = 8'hC;
                    16'hC04D: data_out = 8'hD;
                    16'hC04E: data_out = 8'hE;
                    16'hC04F: data_out = 8'hF;
                    16'hC050: data_out = 8'h10;
                    16'hC051: data_out = 8'h11;
                    16'hC052: data_out = 8'h12;
                    16'hC053: data_out = 8'h13;
                    16'hC054: data_out = 8'h14;
                    16'hC055: data_out = 8'h15;
                    16'hC056: data_out = 8'h16;
                    16'hC057: data_out = 8'h17;
                    16'hC058: data_out = 8'h18;
                    16'hC059: data_out = 8'h19;
                    16'hC05A: data_out = 8'h1A;
                    16'hC05B: data_out = 8'h1B;
                    16'hC05C: data_out = 8'h1C;
                    16'hC05D: data_out = 8'h1D;
                    16'hC05E: data_out = 8'h1E;
                    16'hC05F: data_out = 8'h1F;
                    16'hC060: data_out = 8'h20;
                    16'hC061: data_out = 8'h21;
                    16'hC062: data_out = 8'h22;
                    16'hC063: data_out = 8'h23;
                    16'hC064: data_out = 8'h24;
                    16'hC065: data_out = 8'h25;
                    16'hC066: data_out = 8'h26;
                    16'hC067: data_out = 8'h27;
                    16'hC068: data_out = 8'h28;
                    16'hC069: data_out = 8'h29;
                    16'hC06A: data_out = 8'h2A;
                    16'hC06B: data_out = 8'h2B;
                    16'hC06C: data_out = 8'h2C;
                    16'hC06D: data_out = 8'h2D;
                    16'hC06E: data_out = 8'h2E;
                    16'hC06F: data_out = 8'h2F;
                    16'hC070: data_out = 8'h30;
                    16'hC071: data_out = 8'h31;
                    16'hC072: data_out = 8'h32;
                    16'hC073: data_out = 8'h33;
                    16'hC074: data_out = 8'h34;
                    16'hC075: data_out = 8'h35;
                    16'hC076: data_out = 8'h36;
                    16'hC077: data_out = 8'h37;
                    16'hC078: data_out = 8'h38;
                    16'hC079: data_out = 8'h39;
                    16'hC07A: data_out = 8'h3A;
                    16'hC07B: data_out = 8'h3B;
                    16'hC07C: data_out = 8'h3C;
                    16'hC07D: data_out = 8'h3D;
                    16'hC07E: data_out = 8'h3E;
                    16'hC07F: data_out = 8'h3F;
                    16'hC080: data_out = 8'hC0;
                    16'hC081: data_out = 8'hC1;
                    16'hC082: data_out = 8'hC2;
                    16'hC083: data_out = 8'hC3;
                    16'hC084: data_out = 8'hC4;
                    16'hC085: data_out = 8'hC5;
                    16'hC086: data_out = 8'hC6;
                    16'hC087: data_out = 8'hC7;
                    16'hC088: data_out = 8'hC8;
                    16'hC089: data_out = 8'hC9;
                    16'hC08A: data_out = 8'hCA;
                    16'hC08B: data_out = 8'hCB;
                    16'hC08C: data_out = 8'hCC;
                    16'hC08D: data_out = 8'hCD;
                    16'hC08E: data_out = 8'hCE;
                    16'hC08F: data_out = 8'hCF;
                    16'hC090: data_out = 8'hD0;
                    16'hC091: data_out = 8'hD1;
                    16'hC092: data_out = 8'hD2;
                    16'hC093: data_out = 8'hD3;
                    16'hC094: data_out = 8'hD4;
                    16'hC095: data_out = 8'hD5;
                    16'hC096: data_out = 8'hD6;
                    16'hC097: data_out = 8'hD7;
                    16'hC098: data_out = 8'hD8;
                    16'hC099: data_out = 8'hD9;
                    16'hC09A: data_out = 8'hDA;
                    16'hC09B: data_out = 8'hDB;
                    16'hC09C: data_out = 8'hDC;
                    16'hC09D: data_out = 8'hDD;
                    16'hC09E: data_out = 8'hDE;
                    16'hC09F: data_out = 8'hDF;
                    16'hC0A0: data_out = 8'hE0;
                    16'hC0A1: data_out = 8'hE1;
                    16'hC0A2: data_out = 8'hE2;
                    16'hC0A3: data_out = 8'hE3;
                    16'hC0A4: data_out = 8'hE4;
                    16'hC0A5: data_out = 8'hE5;
                    16'hC0A6: data_out = 8'hE6;
                    16'hC0A7: data_out = 8'hE7;
                    16'hC0A8: data_out = 8'hE8;
                    16'hC0A9: data_out = 8'hE9;
                    16'hC0AA: data_out = 8'hEA;
                    16'hC0AB: data_out = 8'hEB;
                    16'hC0AC: data_out = 8'hEC;
                    16'hC0AD: data_out = 8'hED;
                    16'hC0AE: data_out = 8'hEE;
                    16'hC0AF: data_out = 8'hEF;
                    16'hC0B0: data_out = 8'hF0;
                    16'hC0B1: data_out = 8'hF1;
                    16'hC0B2: data_out = 8'hF2;
                    16'hC0B3: data_out = 8'hF3;
                    16'hC0B4: data_out = 8'hF4;
                    16'hC0B5: data_out = 8'hF5;
                    16'hC0B6: data_out = 8'hF6;
                    16'hC0B7: data_out = 8'hF7;
                    16'hC0B8: data_out = 8'hF8;
                    16'hC0B9: data_out = 8'hF9;
                    16'hC0BA: data_out = 8'hFA;
                    16'hC0BB: data_out = 8'hFB;
                    16'hC0BC: data_out = 8'hFC;
                    16'hC0BD: data_out = 8'hFD;
                    16'hC0BE: data_out = 8'hFE;
                    16'hC0BF: data_out = 8'hFF;
                    16'hC0C0: data_out = 8'h80;
                    16'hC0C1: data_out = 8'h81;
                    16'hC0C2: data_out = 8'h82;
                    16'hC0C3: data_out = 8'h83;
                    16'hC0C4: data_out = 8'h84;
                    16'hC0C5: data_out = 8'h85;
                    16'hC0C6: data_out = 8'h86;
                    16'hC0C7: data_out = 8'h87;
                    16'hC0C8: data_out = 8'h88;
                    16'hC0C9: data_out = 8'h89;
                    16'hC0CA: data_out = 8'h8A;
                    16'hC0CB: data_out = 8'h8B;
                    16'hC0CC: data_out = 8'h8C;
                    16'hC0CD: data_out = 8'h8D;
                    16'hC0CE: data_out = 8'h8E;
                    16'hC0CF: data_out = 8'h8F;
                    16'hC0D0: data_out = 8'h90;
                    16'hC0D1: data_out = 8'h91;
                    16'hC0D2: data_out = 8'h92;
                    16'hC0D3: data_out = 8'h93;
                    16'hC0D4: data_out = 8'h94;
                    16'hC0D5: data_out = 8'h95;
                    16'hC0D6: data_out = 8'h96;
                    16'hC0D7: data_out = 8'h97;
                    16'hC0D8: data_out = 8'h98;
                    16'hC0D9: data_out = 8'h99;
                    16'hC0DA: data_out = 8'h9A;
                    16'hC0DB: data_out = 8'h9B;
                    16'hC0DC: data_out = 8'h9C;
                    16'hC0DD: data_out = 8'h9D;
                    16'hC0DE: data_out = 8'h9E;
                    16'hC0DF: data_out = 8'h9F;
                    16'hC0E0: data_out = 8'hA0;
                    16'hC0E1: data_out = 8'hA1;
                    16'hC0E2: data_out = 8'hA2;
                    16'hC0E3: data_out = 8'hA3;
                    16'hC0E4: data_out = 8'hA4;
                    16'hC0E5: data_out = 8'hA5;
                    16'hC0E6: data_out = 8'hA6;
                    16'hC0E7: data_out = 8'hA7;
                    16'hC0E8: data_out = 8'hA8;
                    16'hC0E9: data_out = 8'hA9;
                    16'hC0EA: data_out = 8'hAA;
                    16'hC0EB: data_out = 8'hAB;
                    16'hC0EC: data_out = 8'hAC;
                    16'hC0ED: data_out = 8'hAD;
                    16'hC0EE: data_out = 8'hAE;
                    16'hC0EF: data_out = 8'hAF;
                    16'hC0F0: data_out = 8'hB0;
                    16'hC0F1: data_out = 8'hB1;
                    16'hC0F2: data_out = 8'hB2;
                    16'hC0F3: data_out = 8'hB3;
                    16'hC0F4: data_out = 8'hB4;
                    16'hC0F5: data_out = 8'hB5;
                    16'hC0F6: data_out = 8'hB6;
                    16'hC0F7: data_out = 8'hB7;
                    16'hC0F8: data_out = 8'hB8;
                    16'hC0F9: data_out = 8'hB9;
                    16'hC0FA: data_out = 8'hBA;
                    16'hC0FB: data_out = 8'hBB;
                    16'hC0FC: data_out = 8'hBC;
                    16'hC0FD: data_out = 8'hBD;
                    16'hC0FE: data_out = 8'hBE;
                    16'hC0FF: data_out = 8'hBF;
                    16'hC100: data_out = 8'hC1;
                    16'hC101: data_out = 8'hC0;
                    16'hC102: data_out = 8'hBF;
                    16'hC103: data_out = 8'hBE;
                    16'hC104: data_out = 8'hBD;
                    16'hC105: data_out = 8'hBC;
                    16'hC106: data_out = 8'hBB;
                    16'hC107: data_out = 8'hBA;
                    16'hC108: data_out = 8'hB9;
                    16'hC109: data_out = 8'hB8;
                    16'hC10A: data_out = 8'hB7;
                    16'hC10B: data_out = 8'hB6;
                    16'hC10C: data_out = 8'hB5;
                    16'hC10D: data_out = 8'hB4;
                    16'hC10E: data_out = 8'hB3;
                    16'hC10F: data_out = 8'hB2;
                    16'hC110: data_out = 8'hB1;
                    16'hC111: data_out = 8'hB0;
                    16'hC112: data_out = 8'hAF;
                    16'hC113: data_out = 8'hAE;
                    16'hC114: data_out = 8'hAD;
                    16'hC115: data_out = 8'hAC;
                    16'hC116: data_out = 8'hAB;
                    16'hC117: data_out = 8'hAA;
                    16'hC118: data_out = 8'hA9;
                    16'hC119: data_out = 8'hA8;
                    16'hC11A: data_out = 8'hA7;
                    16'hC11B: data_out = 8'hA6;
                    16'hC11C: data_out = 8'hA5;
                    16'hC11D: data_out = 8'hA4;
                    16'hC11E: data_out = 8'hA3;
                    16'hC11F: data_out = 8'hA2;
                    16'hC120: data_out = 8'hA1;
                    16'hC121: data_out = 8'hA0;
                    16'hC122: data_out = 8'h9F;
                    16'hC123: data_out = 8'h9E;
                    16'hC124: data_out = 8'h9D;
                    16'hC125: data_out = 8'h9C;
                    16'hC126: data_out = 8'h9B;
                    16'hC127: data_out = 8'h9A;
                    16'hC128: data_out = 8'h99;
                    16'hC129: data_out = 8'h98;
                    16'hC12A: data_out = 8'h97;
                    16'hC12B: data_out = 8'h96;
                    16'hC12C: data_out = 8'h95;
                    16'hC12D: data_out = 8'h94;
                    16'hC12E: data_out = 8'h93;
                    16'hC12F: data_out = 8'h92;
                    16'hC130: data_out = 8'h91;
                    16'hC131: data_out = 8'h90;
                    16'hC132: data_out = 8'h8F;
                    16'hC133: data_out = 8'h8E;
                    16'hC134: data_out = 8'h8D;
                    16'hC135: data_out = 8'h8C;
                    16'hC136: data_out = 8'h8B;
                    16'hC137: data_out = 8'h8A;
                    16'hC138: data_out = 8'h89;
                    16'hC139: data_out = 8'h88;
                    16'hC13A: data_out = 8'h87;
                    16'hC13B: data_out = 8'h86;
                    16'hC13C: data_out = 8'h85;
                    16'hC13D: data_out = 8'h84;
                    16'hC13E: data_out = 8'h83;
                    16'hC13F: data_out = 8'h82;
                    16'hC140: data_out = 8'h81;
                    16'hC141: data_out = 8'h0;
                    16'hC142: data_out = 8'h1;
                    16'hC143: data_out = 8'h2;
                    16'hC144: data_out = 8'h3;
                    16'hC145: data_out = 8'h4;
                    16'hC146: data_out = 8'h5;
                    16'hC147: data_out = 8'h6;
                    16'hC148: data_out = 8'h7;
                    16'hC149: data_out = 8'h8;
                    16'hC14A: data_out = 8'h9;
                    16'hC14B: data_out = 8'hA;
                    16'hC14C: data_out = 8'hB;
                    16'hC14D: data_out = 8'hC;
                    16'hC14E: data_out = 8'hD;
                    16'hC14F: data_out = 8'hE;
                    16'hC150: data_out = 8'hF;
                    16'hC151: data_out = 8'h10;
                    16'hC152: data_out = 8'h11;
                    16'hC153: data_out = 8'h12;
                    16'hC154: data_out = 8'h13;
                    16'hC155: data_out = 8'h14;
                    16'hC156: data_out = 8'h15;
                    16'hC157: data_out = 8'h16;
                    16'hC158: data_out = 8'h17;
                    16'hC159: data_out = 8'h18;
                    16'hC15A: data_out = 8'h19;
                    16'hC15B: data_out = 8'h1A;
                    16'hC15C: data_out = 8'h1B;
                    16'hC15D: data_out = 8'h1C;
                    16'hC15E: data_out = 8'h1D;
                    16'hC15F: data_out = 8'h1E;
                    16'hC160: data_out = 8'h1F;
                    16'hC161: data_out = 8'h20;
                    16'hC162: data_out = 8'h21;
                    16'hC163: data_out = 8'h22;
                    16'hC164: data_out = 8'h23;
                    16'hC165: data_out = 8'h24;
                    16'hC166: data_out = 8'h25;
                    16'hC167: data_out = 8'h26;
                    16'hC168: data_out = 8'h27;
                    16'hC169: data_out = 8'h28;
                    16'hC16A: data_out = 8'h29;
                    16'hC16B: data_out = 8'h2A;
                    16'hC16C: data_out = 8'h2B;
                    16'hC16D: data_out = 8'h2C;
                    16'hC16E: data_out = 8'h2D;
                    16'hC16F: data_out = 8'h2E;
                    16'hC170: data_out = 8'h2F;
                    16'hC171: data_out = 8'h30;
                    16'hC172: data_out = 8'h31;
                    16'hC173: data_out = 8'h32;
                    16'hC174: data_out = 8'h33;
                    16'hC175: data_out = 8'h34;
                    16'hC176: data_out = 8'h35;
                    16'hC177: data_out = 8'h36;
                    16'hC178: data_out = 8'h37;
                    16'hC179: data_out = 8'h38;
                    16'hC17A: data_out = 8'h39;
                    16'hC17B: data_out = 8'h3A;
                    16'hC17C: data_out = 8'h3B;
                    16'hC17D: data_out = 8'h3C;
                    16'hC17E: data_out = 8'h3D;
                    16'hC17F: data_out = 8'h3E;
                    16'hC180: data_out = 8'hC1;
                    16'hC181: data_out = 8'hC2;
                    16'hC182: data_out = 8'hC3;
                    16'hC183: data_out = 8'hC4;
                    16'hC184: data_out = 8'hC5;
                    16'hC185: data_out = 8'hC6;
                    16'hC186: data_out = 8'hC7;
                    16'hC187: data_out = 8'hC8;
                    16'hC188: data_out = 8'hC9;
                    16'hC189: data_out = 8'hCA;
                    16'hC18A: data_out = 8'hCB;
                    16'hC18B: data_out = 8'hCC;
                    16'hC18C: data_out = 8'hCD;
                    16'hC18D: data_out = 8'hCE;
                    16'hC18E: data_out = 8'hCF;
                    16'hC18F: data_out = 8'hD0;
                    16'hC190: data_out = 8'hD1;
                    16'hC191: data_out = 8'hD2;
                    16'hC192: data_out = 8'hD3;
                    16'hC193: data_out = 8'hD4;
                    16'hC194: data_out = 8'hD5;
                    16'hC195: data_out = 8'hD6;
                    16'hC196: data_out = 8'hD7;
                    16'hC197: data_out = 8'hD8;
                    16'hC198: data_out = 8'hD9;
                    16'hC199: data_out = 8'hDA;
                    16'hC19A: data_out = 8'hDB;
                    16'hC19B: data_out = 8'hDC;
                    16'hC19C: data_out = 8'hDD;
                    16'hC19D: data_out = 8'hDE;
                    16'hC19E: data_out = 8'hDF;
                    16'hC19F: data_out = 8'hE0;
                    16'hC1A0: data_out = 8'hE1;
                    16'hC1A1: data_out = 8'hE2;
                    16'hC1A2: data_out = 8'hE3;
                    16'hC1A3: data_out = 8'hE4;
                    16'hC1A4: data_out = 8'hE5;
                    16'hC1A5: data_out = 8'hE6;
                    16'hC1A6: data_out = 8'hE7;
                    16'hC1A7: data_out = 8'hE8;
                    16'hC1A8: data_out = 8'hE9;
                    16'hC1A9: data_out = 8'hEA;
                    16'hC1AA: data_out = 8'hEB;
                    16'hC1AB: data_out = 8'hEC;
                    16'hC1AC: data_out = 8'hED;
                    16'hC1AD: data_out = 8'hEE;
                    16'hC1AE: data_out = 8'hEF;
                    16'hC1AF: data_out = 8'hF0;
                    16'hC1B0: data_out = 8'hF1;
                    16'hC1B1: data_out = 8'hF2;
                    16'hC1B2: data_out = 8'hF3;
                    16'hC1B3: data_out = 8'hF4;
                    16'hC1B4: data_out = 8'hF5;
                    16'hC1B5: data_out = 8'hF6;
                    16'hC1B6: data_out = 8'hF7;
                    16'hC1B7: data_out = 8'hF8;
                    16'hC1B8: data_out = 8'hF9;
                    16'hC1B9: data_out = 8'hFA;
                    16'hC1BA: data_out = 8'hFB;
                    16'hC1BB: data_out = 8'hFC;
                    16'hC1BC: data_out = 8'hFD;
                    16'hC1BD: data_out = 8'hFE;
                    16'hC1BE: data_out = 8'hFF;
                    16'hC1BF: data_out = 8'h80;
                    16'hC1C0: data_out = 8'h81;
                    16'hC1C1: data_out = 8'h82;
                    16'hC1C2: data_out = 8'h83;
                    16'hC1C3: data_out = 8'h84;
                    16'hC1C4: data_out = 8'h85;
                    16'hC1C5: data_out = 8'h86;
                    16'hC1C6: data_out = 8'h87;
                    16'hC1C7: data_out = 8'h88;
                    16'hC1C8: data_out = 8'h89;
                    16'hC1C9: data_out = 8'h8A;
                    16'hC1CA: data_out = 8'h8B;
                    16'hC1CB: data_out = 8'h8C;
                    16'hC1CC: data_out = 8'h8D;
                    16'hC1CD: data_out = 8'h8E;
                    16'hC1CE: data_out = 8'h8F;
                    16'hC1CF: data_out = 8'h90;
                    16'hC1D0: data_out = 8'h91;
                    16'hC1D1: data_out = 8'h92;
                    16'hC1D2: data_out = 8'h93;
                    16'hC1D3: data_out = 8'h94;
                    16'hC1D4: data_out = 8'h95;
                    16'hC1D5: data_out = 8'h96;
                    16'hC1D6: data_out = 8'h97;
                    16'hC1D7: data_out = 8'h98;
                    16'hC1D8: data_out = 8'h99;
                    16'hC1D9: data_out = 8'h9A;
                    16'hC1DA: data_out = 8'h9B;
                    16'hC1DB: data_out = 8'h9C;
                    16'hC1DC: data_out = 8'h9D;
                    16'hC1DD: data_out = 8'h9E;
                    16'hC1DE: data_out = 8'h9F;
                    16'hC1DF: data_out = 8'hA0;
                    16'hC1E0: data_out = 8'hA1;
                    16'hC1E1: data_out = 8'hA2;
                    16'hC1E2: data_out = 8'hA3;
                    16'hC1E3: data_out = 8'hA4;
                    16'hC1E4: data_out = 8'hA5;
                    16'hC1E5: data_out = 8'hA6;
                    16'hC1E6: data_out = 8'hA7;
                    16'hC1E7: data_out = 8'hA8;
                    16'hC1E8: data_out = 8'hA9;
                    16'hC1E9: data_out = 8'hAA;
                    16'hC1EA: data_out = 8'hAB;
                    16'hC1EB: data_out = 8'hAC;
                    16'hC1EC: data_out = 8'hAD;
                    16'hC1ED: data_out = 8'hAE;
                    16'hC1EE: data_out = 8'hAF;
                    16'hC1EF: data_out = 8'hB0;
                    16'hC1F0: data_out = 8'hB1;
                    16'hC1F1: data_out = 8'hB2;
                    16'hC1F2: data_out = 8'hB3;
                    16'hC1F3: data_out = 8'hB4;
                    16'hC1F4: data_out = 8'hB5;
                    16'hC1F5: data_out = 8'hB6;
                    16'hC1F6: data_out = 8'hB7;
                    16'hC1F7: data_out = 8'hB8;
                    16'hC1F8: data_out = 8'hB9;
                    16'hC1F9: data_out = 8'hBA;
                    16'hC1FA: data_out = 8'hBB;
                    16'hC1FB: data_out = 8'hBC;
                    16'hC1FC: data_out = 8'hBD;
                    16'hC1FD: data_out = 8'hBE;
                    16'hC1FE: data_out = 8'hBF;
                    16'hC1FF: data_out = 8'hC0;
                    16'hC200: data_out = 8'hC2;
                    16'hC201: data_out = 8'hC1;
                    16'hC202: data_out = 8'hC0;
                    16'hC203: data_out = 8'hBF;
                    16'hC204: data_out = 8'hBE;
                    16'hC205: data_out = 8'hBD;
                    16'hC206: data_out = 8'hBC;
                    16'hC207: data_out = 8'hBB;
                    16'hC208: data_out = 8'hBA;
                    16'hC209: data_out = 8'hB9;
                    16'hC20A: data_out = 8'hB8;
                    16'hC20B: data_out = 8'hB7;
                    16'hC20C: data_out = 8'hB6;
                    16'hC20D: data_out = 8'hB5;
                    16'hC20E: data_out = 8'hB4;
                    16'hC20F: data_out = 8'hB3;
                    16'hC210: data_out = 8'hB2;
                    16'hC211: data_out = 8'hB1;
                    16'hC212: data_out = 8'hB0;
                    16'hC213: data_out = 8'hAF;
                    16'hC214: data_out = 8'hAE;
                    16'hC215: data_out = 8'hAD;
                    16'hC216: data_out = 8'hAC;
                    16'hC217: data_out = 8'hAB;
                    16'hC218: data_out = 8'hAA;
                    16'hC219: data_out = 8'hA9;
                    16'hC21A: data_out = 8'hA8;
                    16'hC21B: data_out = 8'hA7;
                    16'hC21C: data_out = 8'hA6;
                    16'hC21D: data_out = 8'hA5;
                    16'hC21E: data_out = 8'hA4;
                    16'hC21F: data_out = 8'hA3;
                    16'hC220: data_out = 8'hA2;
                    16'hC221: data_out = 8'hA1;
                    16'hC222: data_out = 8'hA0;
                    16'hC223: data_out = 8'h9F;
                    16'hC224: data_out = 8'h9E;
                    16'hC225: data_out = 8'h9D;
                    16'hC226: data_out = 8'h9C;
                    16'hC227: data_out = 8'h9B;
                    16'hC228: data_out = 8'h9A;
                    16'hC229: data_out = 8'h99;
                    16'hC22A: data_out = 8'h98;
                    16'hC22B: data_out = 8'h97;
                    16'hC22C: data_out = 8'h96;
                    16'hC22D: data_out = 8'h95;
                    16'hC22E: data_out = 8'h94;
                    16'hC22F: data_out = 8'h93;
                    16'hC230: data_out = 8'h92;
                    16'hC231: data_out = 8'h91;
                    16'hC232: data_out = 8'h90;
                    16'hC233: data_out = 8'h8F;
                    16'hC234: data_out = 8'h8E;
                    16'hC235: data_out = 8'h8D;
                    16'hC236: data_out = 8'h8C;
                    16'hC237: data_out = 8'h8B;
                    16'hC238: data_out = 8'h8A;
                    16'hC239: data_out = 8'h89;
                    16'hC23A: data_out = 8'h88;
                    16'hC23B: data_out = 8'h87;
                    16'hC23C: data_out = 8'h86;
                    16'hC23D: data_out = 8'h85;
                    16'hC23E: data_out = 8'h84;
                    16'hC23F: data_out = 8'h83;
                    16'hC240: data_out = 8'h82;
                    16'hC241: data_out = 8'h81;
                    16'hC242: data_out = 8'h0;
                    16'hC243: data_out = 8'h1;
                    16'hC244: data_out = 8'h2;
                    16'hC245: data_out = 8'h3;
                    16'hC246: data_out = 8'h4;
                    16'hC247: data_out = 8'h5;
                    16'hC248: data_out = 8'h6;
                    16'hC249: data_out = 8'h7;
                    16'hC24A: data_out = 8'h8;
                    16'hC24B: data_out = 8'h9;
                    16'hC24C: data_out = 8'hA;
                    16'hC24D: data_out = 8'hB;
                    16'hC24E: data_out = 8'hC;
                    16'hC24F: data_out = 8'hD;
                    16'hC250: data_out = 8'hE;
                    16'hC251: data_out = 8'hF;
                    16'hC252: data_out = 8'h10;
                    16'hC253: data_out = 8'h11;
                    16'hC254: data_out = 8'h12;
                    16'hC255: data_out = 8'h13;
                    16'hC256: data_out = 8'h14;
                    16'hC257: data_out = 8'h15;
                    16'hC258: data_out = 8'h16;
                    16'hC259: data_out = 8'h17;
                    16'hC25A: data_out = 8'h18;
                    16'hC25B: data_out = 8'h19;
                    16'hC25C: data_out = 8'h1A;
                    16'hC25D: data_out = 8'h1B;
                    16'hC25E: data_out = 8'h1C;
                    16'hC25F: data_out = 8'h1D;
                    16'hC260: data_out = 8'h1E;
                    16'hC261: data_out = 8'h1F;
                    16'hC262: data_out = 8'h20;
                    16'hC263: data_out = 8'h21;
                    16'hC264: data_out = 8'h22;
                    16'hC265: data_out = 8'h23;
                    16'hC266: data_out = 8'h24;
                    16'hC267: data_out = 8'h25;
                    16'hC268: data_out = 8'h26;
                    16'hC269: data_out = 8'h27;
                    16'hC26A: data_out = 8'h28;
                    16'hC26B: data_out = 8'h29;
                    16'hC26C: data_out = 8'h2A;
                    16'hC26D: data_out = 8'h2B;
                    16'hC26E: data_out = 8'h2C;
                    16'hC26F: data_out = 8'h2D;
                    16'hC270: data_out = 8'h2E;
                    16'hC271: data_out = 8'h2F;
                    16'hC272: data_out = 8'h30;
                    16'hC273: data_out = 8'h31;
                    16'hC274: data_out = 8'h32;
                    16'hC275: data_out = 8'h33;
                    16'hC276: data_out = 8'h34;
                    16'hC277: data_out = 8'h35;
                    16'hC278: data_out = 8'h36;
                    16'hC279: data_out = 8'h37;
                    16'hC27A: data_out = 8'h38;
                    16'hC27B: data_out = 8'h39;
                    16'hC27C: data_out = 8'h3A;
                    16'hC27D: data_out = 8'h3B;
                    16'hC27E: data_out = 8'h3C;
                    16'hC27F: data_out = 8'h3D;
                    16'hC280: data_out = 8'hC2;
                    16'hC281: data_out = 8'hC3;
                    16'hC282: data_out = 8'hC4;
                    16'hC283: data_out = 8'hC5;
                    16'hC284: data_out = 8'hC6;
                    16'hC285: data_out = 8'hC7;
                    16'hC286: data_out = 8'hC8;
                    16'hC287: data_out = 8'hC9;
                    16'hC288: data_out = 8'hCA;
                    16'hC289: data_out = 8'hCB;
                    16'hC28A: data_out = 8'hCC;
                    16'hC28B: data_out = 8'hCD;
                    16'hC28C: data_out = 8'hCE;
                    16'hC28D: data_out = 8'hCF;
                    16'hC28E: data_out = 8'hD0;
                    16'hC28F: data_out = 8'hD1;
                    16'hC290: data_out = 8'hD2;
                    16'hC291: data_out = 8'hD3;
                    16'hC292: data_out = 8'hD4;
                    16'hC293: data_out = 8'hD5;
                    16'hC294: data_out = 8'hD6;
                    16'hC295: data_out = 8'hD7;
                    16'hC296: data_out = 8'hD8;
                    16'hC297: data_out = 8'hD9;
                    16'hC298: data_out = 8'hDA;
                    16'hC299: data_out = 8'hDB;
                    16'hC29A: data_out = 8'hDC;
                    16'hC29B: data_out = 8'hDD;
                    16'hC29C: data_out = 8'hDE;
                    16'hC29D: data_out = 8'hDF;
                    16'hC29E: data_out = 8'hE0;
                    16'hC29F: data_out = 8'hE1;
                    16'hC2A0: data_out = 8'hE2;
                    16'hC2A1: data_out = 8'hE3;
                    16'hC2A2: data_out = 8'hE4;
                    16'hC2A3: data_out = 8'hE5;
                    16'hC2A4: data_out = 8'hE6;
                    16'hC2A5: data_out = 8'hE7;
                    16'hC2A6: data_out = 8'hE8;
                    16'hC2A7: data_out = 8'hE9;
                    16'hC2A8: data_out = 8'hEA;
                    16'hC2A9: data_out = 8'hEB;
                    16'hC2AA: data_out = 8'hEC;
                    16'hC2AB: data_out = 8'hED;
                    16'hC2AC: data_out = 8'hEE;
                    16'hC2AD: data_out = 8'hEF;
                    16'hC2AE: data_out = 8'hF0;
                    16'hC2AF: data_out = 8'hF1;
                    16'hC2B0: data_out = 8'hF2;
                    16'hC2B1: data_out = 8'hF3;
                    16'hC2B2: data_out = 8'hF4;
                    16'hC2B3: data_out = 8'hF5;
                    16'hC2B4: data_out = 8'hF6;
                    16'hC2B5: data_out = 8'hF7;
                    16'hC2B6: data_out = 8'hF8;
                    16'hC2B7: data_out = 8'hF9;
                    16'hC2B8: data_out = 8'hFA;
                    16'hC2B9: data_out = 8'hFB;
                    16'hC2BA: data_out = 8'hFC;
                    16'hC2BB: data_out = 8'hFD;
                    16'hC2BC: data_out = 8'hFE;
                    16'hC2BD: data_out = 8'hFF;
                    16'hC2BE: data_out = 8'h80;
                    16'hC2BF: data_out = 8'h81;
                    16'hC2C0: data_out = 8'h82;
                    16'hC2C1: data_out = 8'h83;
                    16'hC2C2: data_out = 8'h84;
                    16'hC2C3: data_out = 8'h85;
                    16'hC2C4: data_out = 8'h86;
                    16'hC2C5: data_out = 8'h87;
                    16'hC2C6: data_out = 8'h88;
                    16'hC2C7: data_out = 8'h89;
                    16'hC2C8: data_out = 8'h8A;
                    16'hC2C9: data_out = 8'h8B;
                    16'hC2CA: data_out = 8'h8C;
                    16'hC2CB: data_out = 8'h8D;
                    16'hC2CC: data_out = 8'h8E;
                    16'hC2CD: data_out = 8'h8F;
                    16'hC2CE: data_out = 8'h90;
                    16'hC2CF: data_out = 8'h91;
                    16'hC2D0: data_out = 8'h92;
                    16'hC2D1: data_out = 8'h93;
                    16'hC2D2: data_out = 8'h94;
                    16'hC2D3: data_out = 8'h95;
                    16'hC2D4: data_out = 8'h96;
                    16'hC2D5: data_out = 8'h97;
                    16'hC2D6: data_out = 8'h98;
                    16'hC2D7: data_out = 8'h99;
                    16'hC2D8: data_out = 8'h9A;
                    16'hC2D9: data_out = 8'h9B;
                    16'hC2DA: data_out = 8'h9C;
                    16'hC2DB: data_out = 8'h9D;
                    16'hC2DC: data_out = 8'h9E;
                    16'hC2DD: data_out = 8'h9F;
                    16'hC2DE: data_out = 8'hA0;
                    16'hC2DF: data_out = 8'hA1;
                    16'hC2E0: data_out = 8'hA2;
                    16'hC2E1: data_out = 8'hA3;
                    16'hC2E2: data_out = 8'hA4;
                    16'hC2E3: data_out = 8'hA5;
                    16'hC2E4: data_out = 8'hA6;
                    16'hC2E5: data_out = 8'hA7;
                    16'hC2E6: data_out = 8'hA8;
                    16'hC2E7: data_out = 8'hA9;
                    16'hC2E8: data_out = 8'hAA;
                    16'hC2E9: data_out = 8'hAB;
                    16'hC2EA: data_out = 8'hAC;
                    16'hC2EB: data_out = 8'hAD;
                    16'hC2EC: data_out = 8'hAE;
                    16'hC2ED: data_out = 8'hAF;
                    16'hC2EE: data_out = 8'hB0;
                    16'hC2EF: data_out = 8'hB1;
                    16'hC2F0: data_out = 8'hB2;
                    16'hC2F1: data_out = 8'hB3;
                    16'hC2F2: data_out = 8'hB4;
                    16'hC2F3: data_out = 8'hB5;
                    16'hC2F4: data_out = 8'hB6;
                    16'hC2F5: data_out = 8'hB7;
                    16'hC2F6: data_out = 8'hB8;
                    16'hC2F7: data_out = 8'hB9;
                    16'hC2F8: data_out = 8'hBA;
                    16'hC2F9: data_out = 8'hBB;
                    16'hC2FA: data_out = 8'hBC;
                    16'hC2FB: data_out = 8'hBD;
                    16'hC2FC: data_out = 8'hBE;
                    16'hC2FD: data_out = 8'hBF;
                    16'hC2FE: data_out = 8'hC0;
                    16'hC2FF: data_out = 8'hC1;
                    16'hC300: data_out = 8'hC3;
                    16'hC301: data_out = 8'hC2;
                    16'hC302: data_out = 8'hC1;
                    16'hC303: data_out = 8'hC0;
                    16'hC304: data_out = 8'hBF;
                    16'hC305: data_out = 8'hBE;
                    16'hC306: data_out = 8'hBD;
                    16'hC307: data_out = 8'hBC;
                    16'hC308: data_out = 8'hBB;
                    16'hC309: data_out = 8'hBA;
                    16'hC30A: data_out = 8'hB9;
                    16'hC30B: data_out = 8'hB8;
                    16'hC30C: data_out = 8'hB7;
                    16'hC30D: data_out = 8'hB6;
                    16'hC30E: data_out = 8'hB5;
                    16'hC30F: data_out = 8'hB4;
                    16'hC310: data_out = 8'hB3;
                    16'hC311: data_out = 8'hB2;
                    16'hC312: data_out = 8'hB1;
                    16'hC313: data_out = 8'hB0;
                    16'hC314: data_out = 8'hAF;
                    16'hC315: data_out = 8'hAE;
                    16'hC316: data_out = 8'hAD;
                    16'hC317: data_out = 8'hAC;
                    16'hC318: data_out = 8'hAB;
                    16'hC319: data_out = 8'hAA;
                    16'hC31A: data_out = 8'hA9;
                    16'hC31B: data_out = 8'hA8;
                    16'hC31C: data_out = 8'hA7;
                    16'hC31D: data_out = 8'hA6;
                    16'hC31E: data_out = 8'hA5;
                    16'hC31F: data_out = 8'hA4;
                    16'hC320: data_out = 8'hA3;
                    16'hC321: data_out = 8'hA2;
                    16'hC322: data_out = 8'hA1;
                    16'hC323: data_out = 8'hA0;
                    16'hC324: data_out = 8'h9F;
                    16'hC325: data_out = 8'h9E;
                    16'hC326: data_out = 8'h9D;
                    16'hC327: data_out = 8'h9C;
                    16'hC328: data_out = 8'h9B;
                    16'hC329: data_out = 8'h9A;
                    16'hC32A: data_out = 8'h99;
                    16'hC32B: data_out = 8'h98;
                    16'hC32C: data_out = 8'h97;
                    16'hC32D: data_out = 8'h96;
                    16'hC32E: data_out = 8'h95;
                    16'hC32F: data_out = 8'h94;
                    16'hC330: data_out = 8'h93;
                    16'hC331: data_out = 8'h92;
                    16'hC332: data_out = 8'h91;
                    16'hC333: data_out = 8'h90;
                    16'hC334: data_out = 8'h8F;
                    16'hC335: data_out = 8'h8E;
                    16'hC336: data_out = 8'h8D;
                    16'hC337: data_out = 8'h8C;
                    16'hC338: data_out = 8'h8B;
                    16'hC339: data_out = 8'h8A;
                    16'hC33A: data_out = 8'h89;
                    16'hC33B: data_out = 8'h88;
                    16'hC33C: data_out = 8'h87;
                    16'hC33D: data_out = 8'h86;
                    16'hC33E: data_out = 8'h85;
                    16'hC33F: data_out = 8'h84;
                    16'hC340: data_out = 8'h83;
                    16'hC341: data_out = 8'h82;
                    16'hC342: data_out = 8'h81;
                    16'hC343: data_out = 8'h0;
                    16'hC344: data_out = 8'h1;
                    16'hC345: data_out = 8'h2;
                    16'hC346: data_out = 8'h3;
                    16'hC347: data_out = 8'h4;
                    16'hC348: data_out = 8'h5;
                    16'hC349: data_out = 8'h6;
                    16'hC34A: data_out = 8'h7;
                    16'hC34B: data_out = 8'h8;
                    16'hC34C: data_out = 8'h9;
                    16'hC34D: data_out = 8'hA;
                    16'hC34E: data_out = 8'hB;
                    16'hC34F: data_out = 8'hC;
                    16'hC350: data_out = 8'hD;
                    16'hC351: data_out = 8'hE;
                    16'hC352: data_out = 8'hF;
                    16'hC353: data_out = 8'h10;
                    16'hC354: data_out = 8'h11;
                    16'hC355: data_out = 8'h12;
                    16'hC356: data_out = 8'h13;
                    16'hC357: data_out = 8'h14;
                    16'hC358: data_out = 8'h15;
                    16'hC359: data_out = 8'h16;
                    16'hC35A: data_out = 8'h17;
                    16'hC35B: data_out = 8'h18;
                    16'hC35C: data_out = 8'h19;
                    16'hC35D: data_out = 8'h1A;
                    16'hC35E: data_out = 8'h1B;
                    16'hC35F: data_out = 8'h1C;
                    16'hC360: data_out = 8'h1D;
                    16'hC361: data_out = 8'h1E;
                    16'hC362: data_out = 8'h1F;
                    16'hC363: data_out = 8'h20;
                    16'hC364: data_out = 8'h21;
                    16'hC365: data_out = 8'h22;
                    16'hC366: data_out = 8'h23;
                    16'hC367: data_out = 8'h24;
                    16'hC368: data_out = 8'h25;
                    16'hC369: data_out = 8'h26;
                    16'hC36A: data_out = 8'h27;
                    16'hC36B: data_out = 8'h28;
                    16'hC36C: data_out = 8'h29;
                    16'hC36D: data_out = 8'h2A;
                    16'hC36E: data_out = 8'h2B;
                    16'hC36F: data_out = 8'h2C;
                    16'hC370: data_out = 8'h2D;
                    16'hC371: data_out = 8'h2E;
                    16'hC372: data_out = 8'h2F;
                    16'hC373: data_out = 8'h30;
                    16'hC374: data_out = 8'h31;
                    16'hC375: data_out = 8'h32;
                    16'hC376: data_out = 8'h33;
                    16'hC377: data_out = 8'h34;
                    16'hC378: data_out = 8'h35;
                    16'hC379: data_out = 8'h36;
                    16'hC37A: data_out = 8'h37;
                    16'hC37B: data_out = 8'h38;
                    16'hC37C: data_out = 8'h39;
                    16'hC37D: data_out = 8'h3A;
                    16'hC37E: data_out = 8'h3B;
                    16'hC37F: data_out = 8'h3C;
                    16'hC380: data_out = 8'hC3;
                    16'hC381: data_out = 8'hC4;
                    16'hC382: data_out = 8'hC5;
                    16'hC383: data_out = 8'hC6;
                    16'hC384: data_out = 8'hC7;
                    16'hC385: data_out = 8'hC8;
                    16'hC386: data_out = 8'hC9;
                    16'hC387: data_out = 8'hCA;
                    16'hC388: data_out = 8'hCB;
                    16'hC389: data_out = 8'hCC;
                    16'hC38A: data_out = 8'hCD;
                    16'hC38B: data_out = 8'hCE;
                    16'hC38C: data_out = 8'hCF;
                    16'hC38D: data_out = 8'hD0;
                    16'hC38E: data_out = 8'hD1;
                    16'hC38F: data_out = 8'hD2;
                    16'hC390: data_out = 8'hD3;
                    16'hC391: data_out = 8'hD4;
                    16'hC392: data_out = 8'hD5;
                    16'hC393: data_out = 8'hD6;
                    16'hC394: data_out = 8'hD7;
                    16'hC395: data_out = 8'hD8;
                    16'hC396: data_out = 8'hD9;
                    16'hC397: data_out = 8'hDA;
                    16'hC398: data_out = 8'hDB;
                    16'hC399: data_out = 8'hDC;
                    16'hC39A: data_out = 8'hDD;
                    16'hC39B: data_out = 8'hDE;
                    16'hC39C: data_out = 8'hDF;
                    16'hC39D: data_out = 8'hE0;
                    16'hC39E: data_out = 8'hE1;
                    16'hC39F: data_out = 8'hE2;
                    16'hC3A0: data_out = 8'hE3;
                    16'hC3A1: data_out = 8'hE4;
                    16'hC3A2: data_out = 8'hE5;
                    16'hC3A3: data_out = 8'hE6;
                    16'hC3A4: data_out = 8'hE7;
                    16'hC3A5: data_out = 8'hE8;
                    16'hC3A6: data_out = 8'hE9;
                    16'hC3A7: data_out = 8'hEA;
                    16'hC3A8: data_out = 8'hEB;
                    16'hC3A9: data_out = 8'hEC;
                    16'hC3AA: data_out = 8'hED;
                    16'hC3AB: data_out = 8'hEE;
                    16'hC3AC: data_out = 8'hEF;
                    16'hC3AD: data_out = 8'hF0;
                    16'hC3AE: data_out = 8'hF1;
                    16'hC3AF: data_out = 8'hF2;
                    16'hC3B0: data_out = 8'hF3;
                    16'hC3B1: data_out = 8'hF4;
                    16'hC3B2: data_out = 8'hF5;
                    16'hC3B3: data_out = 8'hF6;
                    16'hC3B4: data_out = 8'hF7;
                    16'hC3B5: data_out = 8'hF8;
                    16'hC3B6: data_out = 8'hF9;
                    16'hC3B7: data_out = 8'hFA;
                    16'hC3B8: data_out = 8'hFB;
                    16'hC3B9: data_out = 8'hFC;
                    16'hC3BA: data_out = 8'hFD;
                    16'hC3BB: data_out = 8'hFE;
                    16'hC3BC: data_out = 8'hFF;
                    16'hC3BD: data_out = 8'h80;
                    16'hC3BE: data_out = 8'h81;
                    16'hC3BF: data_out = 8'h82;
                    16'hC3C0: data_out = 8'h83;
                    16'hC3C1: data_out = 8'h84;
                    16'hC3C2: data_out = 8'h85;
                    16'hC3C3: data_out = 8'h86;
                    16'hC3C4: data_out = 8'h87;
                    16'hC3C5: data_out = 8'h88;
                    16'hC3C6: data_out = 8'h89;
                    16'hC3C7: data_out = 8'h8A;
                    16'hC3C8: data_out = 8'h8B;
                    16'hC3C9: data_out = 8'h8C;
                    16'hC3CA: data_out = 8'h8D;
                    16'hC3CB: data_out = 8'h8E;
                    16'hC3CC: data_out = 8'h8F;
                    16'hC3CD: data_out = 8'h90;
                    16'hC3CE: data_out = 8'h91;
                    16'hC3CF: data_out = 8'h92;
                    16'hC3D0: data_out = 8'h93;
                    16'hC3D1: data_out = 8'h94;
                    16'hC3D2: data_out = 8'h95;
                    16'hC3D3: data_out = 8'h96;
                    16'hC3D4: data_out = 8'h97;
                    16'hC3D5: data_out = 8'h98;
                    16'hC3D6: data_out = 8'h99;
                    16'hC3D7: data_out = 8'h9A;
                    16'hC3D8: data_out = 8'h9B;
                    16'hC3D9: data_out = 8'h9C;
                    16'hC3DA: data_out = 8'h9D;
                    16'hC3DB: data_out = 8'h9E;
                    16'hC3DC: data_out = 8'h9F;
                    16'hC3DD: data_out = 8'hA0;
                    16'hC3DE: data_out = 8'hA1;
                    16'hC3DF: data_out = 8'hA2;
                    16'hC3E0: data_out = 8'hA3;
                    16'hC3E1: data_out = 8'hA4;
                    16'hC3E2: data_out = 8'hA5;
                    16'hC3E3: data_out = 8'hA6;
                    16'hC3E4: data_out = 8'hA7;
                    16'hC3E5: data_out = 8'hA8;
                    16'hC3E6: data_out = 8'hA9;
                    16'hC3E7: data_out = 8'hAA;
                    16'hC3E8: data_out = 8'hAB;
                    16'hC3E9: data_out = 8'hAC;
                    16'hC3EA: data_out = 8'hAD;
                    16'hC3EB: data_out = 8'hAE;
                    16'hC3EC: data_out = 8'hAF;
                    16'hC3ED: data_out = 8'hB0;
                    16'hC3EE: data_out = 8'hB1;
                    16'hC3EF: data_out = 8'hB2;
                    16'hC3F0: data_out = 8'hB3;
                    16'hC3F1: data_out = 8'hB4;
                    16'hC3F2: data_out = 8'hB5;
                    16'hC3F3: data_out = 8'hB6;
                    16'hC3F4: data_out = 8'hB7;
                    16'hC3F5: data_out = 8'hB8;
                    16'hC3F6: data_out = 8'hB9;
                    16'hC3F7: data_out = 8'hBA;
                    16'hC3F8: data_out = 8'hBB;
                    16'hC3F9: data_out = 8'hBC;
                    16'hC3FA: data_out = 8'hBD;
                    16'hC3FB: data_out = 8'hBE;
                    16'hC3FC: data_out = 8'hBF;
                    16'hC3FD: data_out = 8'hC0;
                    16'hC3FE: data_out = 8'hC1;
                    16'hC3FF: data_out = 8'hC2;
                    16'hC400: data_out = 8'hC4;
                    16'hC401: data_out = 8'hC3;
                    16'hC402: data_out = 8'hC2;
                    16'hC403: data_out = 8'hC1;
                    16'hC404: data_out = 8'hC0;
                    16'hC405: data_out = 8'hBF;
                    16'hC406: data_out = 8'hBE;
                    16'hC407: data_out = 8'hBD;
                    16'hC408: data_out = 8'hBC;
                    16'hC409: data_out = 8'hBB;
                    16'hC40A: data_out = 8'hBA;
                    16'hC40B: data_out = 8'hB9;
                    16'hC40C: data_out = 8'hB8;
                    16'hC40D: data_out = 8'hB7;
                    16'hC40E: data_out = 8'hB6;
                    16'hC40F: data_out = 8'hB5;
                    16'hC410: data_out = 8'hB4;
                    16'hC411: data_out = 8'hB3;
                    16'hC412: data_out = 8'hB2;
                    16'hC413: data_out = 8'hB1;
                    16'hC414: data_out = 8'hB0;
                    16'hC415: data_out = 8'hAF;
                    16'hC416: data_out = 8'hAE;
                    16'hC417: data_out = 8'hAD;
                    16'hC418: data_out = 8'hAC;
                    16'hC419: data_out = 8'hAB;
                    16'hC41A: data_out = 8'hAA;
                    16'hC41B: data_out = 8'hA9;
                    16'hC41C: data_out = 8'hA8;
                    16'hC41D: data_out = 8'hA7;
                    16'hC41E: data_out = 8'hA6;
                    16'hC41F: data_out = 8'hA5;
                    16'hC420: data_out = 8'hA4;
                    16'hC421: data_out = 8'hA3;
                    16'hC422: data_out = 8'hA2;
                    16'hC423: data_out = 8'hA1;
                    16'hC424: data_out = 8'hA0;
                    16'hC425: data_out = 8'h9F;
                    16'hC426: data_out = 8'h9E;
                    16'hC427: data_out = 8'h9D;
                    16'hC428: data_out = 8'h9C;
                    16'hC429: data_out = 8'h9B;
                    16'hC42A: data_out = 8'h9A;
                    16'hC42B: data_out = 8'h99;
                    16'hC42C: data_out = 8'h98;
                    16'hC42D: data_out = 8'h97;
                    16'hC42E: data_out = 8'h96;
                    16'hC42F: data_out = 8'h95;
                    16'hC430: data_out = 8'h94;
                    16'hC431: data_out = 8'h93;
                    16'hC432: data_out = 8'h92;
                    16'hC433: data_out = 8'h91;
                    16'hC434: data_out = 8'h90;
                    16'hC435: data_out = 8'h8F;
                    16'hC436: data_out = 8'h8E;
                    16'hC437: data_out = 8'h8D;
                    16'hC438: data_out = 8'h8C;
                    16'hC439: data_out = 8'h8B;
                    16'hC43A: data_out = 8'h8A;
                    16'hC43B: data_out = 8'h89;
                    16'hC43C: data_out = 8'h88;
                    16'hC43D: data_out = 8'h87;
                    16'hC43E: data_out = 8'h86;
                    16'hC43F: data_out = 8'h85;
                    16'hC440: data_out = 8'h84;
                    16'hC441: data_out = 8'h83;
                    16'hC442: data_out = 8'h82;
                    16'hC443: data_out = 8'h81;
                    16'hC444: data_out = 8'h0;
                    16'hC445: data_out = 8'h1;
                    16'hC446: data_out = 8'h2;
                    16'hC447: data_out = 8'h3;
                    16'hC448: data_out = 8'h4;
                    16'hC449: data_out = 8'h5;
                    16'hC44A: data_out = 8'h6;
                    16'hC44B: data_out = 8'h7;
                    16'hC44C: data_out = 8'h8;
                    16'hC44D: data_out = 8'h9;
                    16'hC44E: data_out = 8'hA;
                    16'hC44F: data_out = 8'hB;
                    16'hC450: data_out = 8'hC;
                    16'hC451: data_out = 8'hD;
                    16'hC452: data_out = 8'hE;
                    16'hC453: data_out = 8'hF;
                    16'hC454: data_out = 8'h10;
                    16'hC455: data_out = 8'h11;
                    16'hC456: data_out = 8'h12;
                    16'hC457: data_out = 8'h13;
                    16'hC458: data_out = 8'h14;
                    16'hC459: data_out = 8'h15;
                    16'hC45A: data_out = 8'h16;
                    16'hC45B: data_out = 8'h17;
                    16'hC45C: data_out = 8'h18;
                    16'hC45D: data_out = 8'h19;
                    16'hC45E: data_out = 8'h1A;
                    16'hC45F: data_out = 8'h1B;
                    16'hC460: data_out = 8'h1C;
                    16'hC461: data_out = 8'h1D;
                    16'hC462: data_out = 8'h1E;
                    16'hC463: data_out = 8'h1F;
                    16'hC464: data_out = 8'h20;
                    16'hC465: data_out = 8'h21;
                    16'hC466: data_out = 8'h22;
                    16'hC467: data_out = 8'h23;
                    16'hC468: data_out = 8'h24;
                    16'hC469: data_out = 8'h25;
                    16'hC46A: data_out = 8'h26;
                    16'hC46B: data_out = 8'h27;
                    16'hC46C: data_out = 8'h28;
                    16'hC46D: data_out = 8'h29;
                    16'hC46E: data_out = 8'h2A;
                    16'hC46F: data_out = 8'h2B;
                    16'hC470: data_out = 8'h2C;
                    16'hC471: data_out = 8'h2D;
                    16'hC472: data_out = 8'h2E;
                    16'hC473: data_out = 8'h2F;
                    16'hC474: data_out = 8'h30;
                    16'hC475: data_out = 8'h31;
                    16'hC476: data_out = 8'h32;
                    16'hC477: data_out = 8'h33;
                    16'hC478: data_out = 8'h34;
                    16'hC479: data_out = 8'h35;
                    16'hC47A: data_out = 8'h36;
                    16'hC47B: data_out = 8'h37;
                    16'hC47C: data_out = 8'h38;
                    16'hC47D: data_out = 8'h39;
                    16'hC47E: data_out = 8'h3A;
                    16'hC47F: data_out = 8'h3B;
                    16'hC480: data_out = 8'hC4;
                    16'hC481: data_out = 8'hC5;
                    16'hC482: data_out = 8'hC6;
                    16'hC483: data_out = 8'hC7;
                    16'hC484: data_out = 8'hC8;
                    16'hC485: data_out = 8'hC9;
                    16'hC486: data_out = 8'hCA;
                    16'hC487: data_out = 8'hCB;
                    16'hC488: data_out = 8'hCC;
                    16'hC489: data_out = 8'hCD;
                    16'hC48A: data_out = 8'hCE;
                    16'hC48B: data_out = 8'hCF;
                    16'hC48C: data_out = 8'hD0;
                    16'hC48D: data_out = 8'hD1;
                    16'hC48E: data_out = 8'hD2;
                    16'hC48F: data_out = 8'hD3;
                    16'hC490: data_out = 8'hD4;
                    16'hC491: data_out = 8'hD5;
                    16'hC492: data_out = 8'hD6;
                    16'hC493: data_out = 8'hD7;
                    16'hC494: data_out = 8'hD8;
                    16'hC495: data_out = 8'hD9;
                    16'hC496: data_out = 8'hDA;
                    16'hC497: data_out = 8'hDB;
                    16'hC498: data_out = 8'hDC;
                    16'hC499: data_out = 8'hDD;
                    16'hC49A: data_out = 8'hDE;
                    16'hC49B: data_out = 8'hDF;
                    16'hC49C: data_out = 8'hE0;
                    16'hC49D: data_out = 8'hE1;
                    16'hC49E: data_out = 8'hE2;
                    16'hC49F: data_out = 8'hE3;
                    16'hC4A0: data_out = 8'hE4;
                    16'hC4A1: data_out = 8'hE5;
                    16'hC4A2: data_out = 8'hE6;
                    16'hC4A3: data_out = 8'hE7;
                    16'hC4A4: data_out = 8'hE8;
                    16'hC4A5: data_out = 8'hE9;
                    16'hC4A6: data_out = 8'hEA;
                    16'hC4A7: data_out = 8'hEB;
                    16'hC4A8: data_out = 8'hEC;
                    16'hC4A9: data_out = 8'hED;
                    16'hC4AA: data_out = 8'hEE;
                    16'hC4AB: data_out = 8'hEF;
                    16'hC4AC: data_out = 8'hF0;
                    16'hC4AD: data_out = 8'hF1;
                    16'hC4AE: data_out = 8'hF2;
                    16'hC4AF: data_out = 8'hF3;
                    16'hC4B0: data_out = 8'hF4;
                    16'hC4B1: data_out = 8'hF5;
                    16'hC4B2: data_out = 8'hF6;
                    16'hC4B3: data_out = 8'hF7;
                    16'hC4B4: data_out = 8'hF8;
                    16'hC4B5: data_out = 8'hF9;
                    16'hC4B6: data_out = 8'hFA;
                    16'hC4B7: data_out = 8'hFB;
                    16'hC4B8: data_out = 8'hFC;
                    16'hC4B9: data_out = 8'hFD;
                    16'hC4BA: data_out = 8'hFE;
                    16'hC4BB: data_out = 8'hFF;
                    16'hC4BC: data_out = 8'h80;
                    16'hC4BD: data_out = 8'h81;
                    16'hC4BE: data_out = 8'h82;
                    16'hC4BF: data_out = 8'h83;
                    16'hC4C0: data_out = 8'h84;
                    16'hC4C1: data_out = 8'h85;
                    16'hC4C2: data_out = 8'h86;
                    16'hC4C3: data_out = 8'h87;
                    16'hC4C4: data_out = 8'h88;
                    16'hC4C5: data_out = 8'h89;
                    16'hC4C6: data_out = 8'h8A;
                    16'hC4C7: data_out = 8'h8B;
                    16'hC4C8: data_out = 8'h8C;
                    16'hC4C9: data_out = 8'h8D;
                    16'hC4CA: data_out = 8'h8E;
                    16'hC4CB: data_out = 8'h8F;
                    16'hC4CC: data_out = 8'h90;
                    16'hC4CD: data_out = 8'h91;
                    16'hC4CE: data_out = 8'h92;
                    16'hC4CF: data_out = 8'h93;
                    16'hC4D0: data_out = 8'h94;
                    16'hC4D1: data_out = 8'h95;
                    16'hC4D2: data_out = 8'h96;
                    16'hC4D3: data_out = 8'h97;
                    16'hC4D4: data_out = 8'h98;
                    16'hC4D5: data_out = 8'h99;
                    16'hC4D6: data_out = 8'h9A;
                    16'hC4D7: data_out = 8'h9B;
                    16'hC4D8: data_out = 8'h9C;
                    16'hC4D9: data_out = 8'h9D;
                    16'hC4DA: data_out = 8'h9E;
                    16'hC4DB: data_out = 8'h9F;
                    16'hC4DC: data_out = 8'hA0;
                    16'hC4DD: data_out = 8'hA1;
                    16'hC4DE: data_out = 8'hA2;
                    16'hC4DF: data_out = 8'hA3;
                    16'hC4E0: data_out = 8'hA4;
                    16'hC4E1: data_out = 8'hA5;
                    16'hC4E2: data_out = 8'hA6;
                    16'hC4E3: data_out = 8'hA7;
                    16'hC4E4: data_out = 8'hA8;
                    16'hC4E5: data_out = 8'hA9;
                    16'hC4E6: data_out = 8'hAA;
                    16'hC4E7: data_out = 8'hAB;
                    16'hC4E8: data_out = 8'hAC;
                    16'hC4E9: data_out = 8'hAD;
                    16'hC4EA: data_out = 8'hAE;
                    16'hC4EB: data_out = 8'hAF;
                    16'hC4EC: data_out = 8'hB0;
                    16'hC4ED: data_out = 8'hB1;
                    16'hC4EE: data_out = 8'hB2;
                    16'hC4EF: data_out = 8'hB3;
                    16'hC4F0: data_out = 8'hB4;
                    16'hC4F1: data_out = 8'hB5;
                    16'hC4F2: data_out = 8'hB6;
                    16'hC4F3: data_out = 8'hB7;
                    16'hC4F4: data_out = 8'hB8;
                    16'hC4F5: data_out = 8'hB9;
                    16'hC4F6: data_out = 8'hBA;
                    16'hC4F7: data_out = 8'hBB;
                    16'hC4F8: data_out = 8'hBC;
                    16'hC4F9: data_out = 8'hBD;
                    16'hC4FA: data_out = 8'hBE;
                    16'hC4FB: data_out = 8'hBF;
                    16'hC4FC: data_out = 8'hC0;
                    16'hC4FD: data_out = 8'hC1;
                    16'hC4FE: data_out = 8'hC2;
                    16'hC4FF: data_out = 8'hC3;
                    16'hC500: data_out = 8'hC5;
                    16'hC501: data_out = 8'hC4;
                    16'hC502: data_out = 8'hC3;
                    16'hC503: data_out = 8'hC2;
                    16'hC504: data_out = 8'hC1;
                    16'hC505: data_out = 8'hC0;
                    16'hC506: data_out = 8'hBF;
                    16'hC507: data_out = 8'hBE;
                    16'hC508: data_out = 8'hBD;
                    16'hC509: data_out = 8'hBC;
                    16'hC50A: data_out = 8'hBB;
                    16'hC50B: data_out = 8'hBA;
                    16'hC50C: data_out = 8'hB9;
                    16'hC50D: data_out = 8'hB8;
                    16'hC50E: data_out = 8'hB7;
                    16'hC50F: data_out = 8'hB6;
                    16'hC510: data_out = 8'hB5;
                    16'hC511: data_out = 8'hB4;
                    16'hC512: data_out = 8'hB3;
                    16'hC513: data_out = 8'hB2;
                    16'hC514: data_out = 8'hB1;
                    16'hC515: data_out = 8'hB0;
                    16'hC516: data_out = 8'hAF;
                    16'hC517: data_out = 8'hAE;
                    16'hC518: data_out = 8'hAD;
                    16'hC519: data_out = 8'hAC;
                    16'hC51A: data_out = 8'hAB;
                    16'hC51B: data_out = 8'hAA;
                    16'hC51C: data_out = 8'hA9;
                    16'hC51D: data_out = 8'hA8;
                    16'hC51E: data_out = 8'hA7;
                    16'hC51F: data_out = 8'hA6;
                    16'hC520: data_out = 8'hA5;
                    16'hC521: data_out = 8'hA4;
                    16'hC522: data_out = 8'hA3;
                    16'hC523: data_out = 8'hA2;
                    16'hC524: data_out = 8'hA1;
                    16'hC525: data_out = 8'hA0;
                    16'hC526: data_out = 8'h9F;
                    16'hC527: data_out = 8'h9E;
                    16'hC528: data_out = 8'h9D;
                    16'hC529: data_out = 8'h9C;
                    16'hC52A: data_out = 8'h9B;
                    16'hC52B: data_out = 8'h9A;
                    16'hC52C: data_out = 8'h99;
                    16'hC52D: data_out = 8'h98;
                    16'hC52E: data_out = 8'h97;
                    16'hC52F: data_out = 8'h96;
                    16'hC530: data_out = 8'h95;
                    16'hC531: data_out = 8'h94;
                    16'hC532: data_out = 8'h93;
                    16'hC533: data_out = 8'h92;
                    16'hC534: data_out = 8'h91;
                    16'hC535: data_out = 8'h90;
                    16'hC536: data_out = 8'h8F;
                    16'hC537: data_out = 8'h8E;
                    16'hC538: data_out = 8'h8D;
                    16'hC539: data_out = 8'h8C;
                    16'hC53A: data_out = 8'h8B;
                    16'hC53B: data_out = 8'h8A;
                    16'hC53C: data_out = 8'h89;
                    16'hC53D: data_out = 8'h88;
                    16'hC53E: data_out = 8'h87;
                    16'hC53F: data_out = 8'h86;
                    16'hC540: data_out = 8'h85;
                    16'hC541: data_out = 8'h84;
                    16'hC542: data_out = 8'h83;
                    16'hC543: data_out = 8'h82;
                    16'hC544: data_out = 8'h81;
                    16'hC545: data_out = 8'h0;
                    16'hC546: data_out = 8'h1;
                    16'hC547: data_out = 8'h2;
                    16'hC548: data_out = 8'h3;
                    16'hC549: data_out = 8'h4;
                    16'hC54A: data_out = 8'h5;
                    16'hC54B: data_out = 8'h6;
                    16'hC54C: data_out = 8'h7;
                    16'hC54D: data_out = 8'h8;
                    16'hC54E: data_out = 8'h9;
                    16'hC54F: data_out = 8'hA;
                    16'hC550: data_out = 8'hB;
                    16'hC551: data_out = 8'hC;
                    16'hC552: data_out = 8'hD;
                    16'hC553: data_out = 8'hE;
                    16'hC554: data_out = 8'hF;
                    16'hC555: data_out = 8'h10;
                    16'hC556: data_out = 8'h11;
                    16'hC557: data_out = 8'h12;
                    16'hC558: data_out = 8'h13;
                    16'hC559: data_out = 8'h14;
                    16'hC55A: data_out = 8'h15;
                    16'hC55B: data_out = 8'h16;
                    16'hC55C: data_out = 8'h17;
                    16'hC55D: data_out = 8'h18;
                    16'hC55E: data_out = 8'h19;
                    16'hC55F: data_out = 8'h1A;
                    16'hC560: data_out = 8'h1B;
                    16'hC561: data_out = 8'h1C;
                    16'hC562: data_out = 8'h1D;
                    16'hC563: data_out = 8'h1E;
                    16'hC564: data_out = 8'h1F;
                    16'hC565: data_out = 8'h20;
                    16'hC566: data_out = 8'h21;
                    16'hC567: data_out = 8'h22;
                    16'hC568: data_out = 8'h23;
                    16'hC569: data_out = 8'h24;
                    16'hC56A: data_out = 8'h25;
                    16'hC56B: data_out = 8'h26;
                    16'hC56C: data_out = 8'h27;
                    16'hC56D: data_out = 8'h28;
                    16'hC56E: data_out = 8'h29;
                    16'hC56F: data_out = 8'h2A;
                    16'hC570: data_out = 8'h2B;
                    16'hC571: data_out = 8'h2C;
                    16'hC572: data_out = 8'h2D;
                    16'hC573: data_out = 8'h2E;
                    16'hC574: data_out = 8'h2F;
                    16'hC575: data_out = 8'h30;
                    16'hC576: data_out = 8'h31;
                    16'hC577: data_out = 8'h32;
                    16'hC578: data_out = 8'h33;
                    16'hC579: data_out = 8'h34;
                    16'hC57A: data_out = 8'h35;
                    16'hC57B: data_out = 8'h36;
                    16'hC57C: data_out = 8'h37;
                    16'hC57D: data_out = 8'h38;
                    16'hC57E: data_out = 8'h39;
                    16'hC57F: data_out = 8'h3A;
                    16'hC580: data_out = 8'hC5;
                    16'hC581: data_out = 8'hC6;
                    16'hC582: data_out = 8'hC7;
                    16'hC583: data_out = 8'hC8;
                    16'hC584: data_out = 8'hC9;
                    16'hC585: data_out = 8'hCA;
                    16'hC586: data_out = 8'hCB;
                    16'hC587: data_out = 8'hCC;
                    16'hC588: data_out = 8'hCD;
                    16'hC589: data_out = 8'hCE;
                    16'hC58A: data_out = 8'hCF;
                    16'hC58B: data_out = 8'hD0;
                    16'hC58C: data_out = 8'hD1;
                    16'hC58D: data_out = 8'hD2;
                    16'hC58E: data_out = 8'hD3;
                    16'hC58F: data_out = 8'hD4;
                    16'hC590: data_out = 8'hD5;
                    16'hC591: data_out = 8'hD6;
                    16'hC592: data_out = 8'hD7;
                    16'hC593: data_out = 8'hD8;
                    16'hC594: data_out = 8'hD9;
                    16'hC595: data_out = 8'hDA;
                    16'hC596: data_out = 8'hDB;
                    16'hC597: data_out = 8'hDC;
                    16'hC598: data_out = 8'hDD;
                    16'hC599: data_out = 8'hDE;
                    16'hC59A: data_out = 8'hDF;
                    16'hC59B: data_out = 8'hE0;
                    16'hC59C: data_out = 8'hE1;
                    16'hC59D: data_out = 8'hE2;
                    16'hC59E: data_out = 8'hE3;
                    16'hC59F: data_out = 8'hE4;
                    16'hC5A0: data_out = 8'hE5;
                    16'hC5A1: data_out = 8'hE6;
                    16'hC5A2: data_out = 8'hE7;
                    16'hC5A3: data_out = 8'hE8;
                    16'hC5A4: data_out = 8'hE9;
                    16'hC5A5: data_out = 8'hEA;
                    16'hC5A6: data_out = 8'hEB;
                    16'hC5A7: data_out = 8'hEC;
                    16'hC5A8: data_out = 8'hED;
                    16'hC5A9: data_out = 8'hEE;
                    16'hC5AA: data_out = 8'hEF;
                    16'hC5AB: data_out = 8'hF0;
                    16'hC5AC: data_out = 8'hF1;
                    16'hC5AD: data_out = 8'hF2;
                    16'hC5AE: data_out = 8'hF3;
                    16'hC5AF: data_out = 8'hF4;
                    16'hC5B0: data_out = 8'hF5;
                    16'hC5B1: data_out = 8'hF6;
                    16'hC5B2: data_out = 8'hF7;
                    16'hC5B3: data_out = 8'hF8;
                    16'hC5B4: data_out = 8'hF9;
                    16'hC5B5: data_out = 8'hFA;
                    16'hC5B6: data_out = 8'hFB;
                    16'hC5B7: data_out = 8'hFC;
                    16'hC5B8: data_out = 8'hFD;
                    16'hC5B9: data_out = 8'hFE;
                    16'hC5BA: data_out = 8'hFF;
                    16'hC5BB: data_out = 8'h80;
                    16'hC5BC: data_out = 8'h81;
                    16'hC5BD: data_out = 8'h82;
                    16'hC5BE: data_out = 8'h83;
                    16'hC5BF: data_out = 8'h84;
                    16'hC5C0: data_out = 8'h85;
                    16'hC5C1: data_out = 8'h86;
                    16'hC5C2: data_out = 8'h87;
                    16'hC5C3: data_out = 8'h88;
                    16'hC5C4: data_out = 8'h89;
                    16'hC5C5: data_out = 8'h8A;
                    16'hC5C6: data_out = 8'h8B;
                    16'hC5C7: data_out = 8'h8C;
                    16'hC5C8: data_out = 8'h8D;
                    16'hC5C9: data_out = 8'h8E;
                    16'hC5CA: data_out = 8'h8F;
                    16'hC5CB: data_out = 8'h90;
                    16'hC5CC: data_out = 8'h91;
                    16'hC5CD: data_out = 8'h92;
                    16'hC5CE: data_out = 8'h93;
                    16'hC5CF: data_out = 8'h94;
                    16'hC5D0: data_out = 8'h95;
                    16'hC5D1: data_out = 8'h96;
                    16'hC5D2: data_out = 8'h97;
                    16'hC5D3: data_out = 8'h98;
                    16'hC5D4: data_out = 8'h99;
                    16'hC5D5: data_out = 8'h9A;
                    16'hC5D6: data_out = 8'h9B;
                    16'hC5D7: data_out = 8'h9C;
                    16'hC5D8: data_out = 8'h9D;
                    16'hC5D9: data_out = 8'h9E;
                    16'hC5DA: data_out = 8'h9F;
                    16'hC5DB: data_out = 8'hA0;
                    16'hC5DC: data_out = 8'hA1;
                    16'hC5DD: data_out = 8'hA2;
                    16'hC5DE: data_out = 8'hA3;
                    16'hC5DF: data_out = 8'hA4;
                    16'hC5E0: data_out = 8'hA5;
                    16'hC5E1: data_out = 8'hA6;
                    16'hC5E2: data_out = 8'hA7;
                    16'hC5E3: data_out = 8'hA8;
                    16'hC5E4: data_out = 8'hA9;
                    16'hC5E5: data_out = 8'hAA;
                    16'hC5E6: data_out = 8'hAB;
                    16'hC5E7: data_out = 8'hAC;
                    16'hC5E8: data_out = 8'hAD;
                    16'hC5E9: data_out = 8'hAE;
                    16'hC5EA: data_out = 8'hAF;
                    16'hC5EB: data_out = 8'hB0;
                    16'hC5EC: data_out = 8'hB1;
                    16'hC5ED: data_out = 8'hB2;
                    16'hC5EE: data_out = 8'hB3;
                    16'hC5EF: data_out = 8'hB4;
                    16'hC5F0: data_out = 8'hB5;
                    16'hC5F1: data_out = 8'hB6;
                    16'hC5F2: data_out = 8'hB7;
                    16'hC5F3: data_out = 8'hB8;
                    16'hC5F4: data_out = 8'hB9;
                    16'hC5F5: data_out = 8'hBA;
                    16'hC5F6: data_out = 8'hBB;
                    16'hC5F7: data_out = 8'hBC;
                    16'hC5F8: data_out = 8'hBD;
                    16'hC5F9: data_out = 8'hBE;
                    16'hC5FA: data_out = 8'hBF;
                    16'hC5FB: data_out = 8'hC0;
                    16'hC5FC: data_out = 8'hC1;
                    16'hC5FD: data_out = 8'hC2;
                    16'hC5FE: data_out = 8'hC3;
                    16'hC5FF: data_out = 8'hC4;
                    16'hC600: data_out = 8'hC6;
                    16'hC601: data_out = 8'hC5;
                    16'hC602: data_out = 8'hC4;
                    16'hC603: data_out = 8'hC3;
                    16'hC604: data_out = 8'hC2;
                    16'hC605: data_out = 8'hC1;
                    16'hC606: data_out = 8'hC0;
                    16'hC607: data_out = 8'hBF;
                    16'hC608: data_out = 8'hBE;
                    16'hC609: data_out = 8'hBD;
                    16'hC60A: data_out = 8'hBC;
                    16'hC60B: data_out = 8'hBB;
                    16'hC60C: data_out = 8'hBA;
                    16'hC60D: data_out = 8'hB9;
                    16'hC60E: data_out = 8'hB8;
                    16'hC60F: data_out = 8'hB7;
                    16'hC610: data_out = 8'hB6;
                    16'hC611: data_out = 8'hB5;
                    16'hC612: data_out = 8'hB4;
                    16'hC613: data_out = 8'hB3;
                    16'hC614: data_out = 8'hB2;
                    16'hC615: data_out = 8'hB1;
                    16'hC616: data_out = 8'hB0;
                    16'hC617: data_out = 8'hAF;
                    16'hC618: data_out = 8'hAE;
                    16'hC619: data_out = 8'hAD;
                    16'hC61A: data_out = 8'hAC;
                    16'hC61B: data_out = 8'hAB;
                    16'hC61C: data_out = 8'hAA;
                    16'hC61D: data_out = 8'hA9;
                    16'hC61E: data_out = 8'hA8;
                    16'hC61F: data_out = 8'hA7;
                    16'hC620: data_out = 8'hA6;
                    16'hC621: data_out = 8'hA5;
                    16'hC622: data_out = 8'hA4;
                    16'hC623: data_out = 8'hA3;
                    16'hC624: data_out = 8'hA2;
                    16'hC625: data_out = 8'hA1;
                    16'hC626: data_out = 8'hA0;
                    16'hC627: data_out = 8'h9F;
                    16'hC628: data_out = 8'h9E;
                    16'hC629: data_out = 8'h9D;
                    16'hC62A: data_out = 8'h9C;
                    16'hC62B: data_out = 8'h9B;
                    16'hC62C: data_out = 8'h9A;
                    16'hC62D: data_out = 8'h99;
                    16'hC62E: data_out = 8'h98;
                    16'hC62F: data_out = 8'h97;
                    16'hC630: data_out = 8'h96;
                    16'hC631: data_out = 8'h95;
                    16'hC632: data_out = 8'h94;
                    16'hC633: data_out = 8'h93;
                    16'hC634: data_out = 8'h92;
                    16'hC635: data_out = 8'h91;
                    16'hC636: data_out = 8'h90;
                    16'hC637: data_out = 8'h8F;
                    16'hC638: data_out = 8'h8E;
                    16'hC639: data_out = 8'h8D;
                    16'hC63A: data_out = 8'h8C;
                    16'hC63B: data_out = 8'h8B;
                    16'hC63C: data_out = 8'h8A;
                    16'hC63D: data_out = 8'h89;
                    16'hC63E: data_out = 8'h88;
                    16'hC63F: data_out = 8'h87;
                    16'hC640: data_out = 8'h86;
                    16'hC641: data_out = 8'h85;
                    16'hC642: data_out = 8'h84;
                    16'hC643: data_out = 8'h83;
                    16'hC644: data_out = 8'h82;
                    16'hC645: data_out = 8'h81;
                    16'hC646: data_out = 8'h0;
                    16'hC647: data_out = 8'h1;
                    16'hC648: data_out = 8'h2;
                    16'hC649: data_out = 8'h3;
                    16'hC64A: data_out = 8'h4;
                    16'hC64B: data_out = 8'h5;
                    16'hC64C: data_out = 8'h6;
                    16'hC64D: data_out = 8'h7;
                    16'hC64E: data_out = 8'h8;
                    16'hC64F: data_out = 8'h9;
                    16'hC650: data_out = 8'hA;
                    16'hC651: data_out = 8'hB;
                    16'hC652: data_out = 8'hC;
                    16'hC653: data_out = 8'hD;
                    16'hC654: data_out = 8'hE;
                    16'hC655: data_out = 8'hF;
                    16'hC656: data_out = 8'h10;
                    16'hC657: data_out = 8'h11;
                    16'hC658: data_out = 8'h12;
                    16'hC659: data_out = 8'h13;
                    16'hC65A: data_out = 8'h14;
                    16'hC65B: data_out = 8'h15;
                    16'hC65C: data_out = 8'h16;
                    16'hC65D: data_out = 8'h17;
                    16'hC65E: data_out = 8'h18;
                    16'hC65F: data_out = 8'h19;
                    16'hC660: data_out = 8'h1A;
                    16'hC661: data_out = 8'h1B;
                    16'hC662: data_out = 8'h1C;
                    16'hC663: data_out = 8'h1D;
                    16'hC664: data_out = 8'h1E;
                    16'hC665: data_out = 8'h1F;
                    16'hC666: data_out = 8'h20;
                    16'hC667: data_out = 8'h21;
                    16'hC668: data_out = 8'h22;
                    16'hC669: data_out = 8'h23;
                    16'hC66A: data_out = 8'h24;
                    16'hC66B: data_out = 8'h25;
                    16'hC66C: data_out = 8'h26;
                    16'hC66D: data_out = 8'h27;
                    16'hC66E: data_out = 8'h28;
                    16'hC66F: data_out = 8'h29;
                    16'hC670: data_out = 8'h2A;
                    16'hC671: data_out = 8'h2B;
                    16'hC672: data_out = 8'h2C;
                    16'hC673: data_out = 8'h2D;
                    16'hC674: data_out = 8'h2E;
                    16'hC675: data_out = 8'h2F;
                    16'hC676: data_out = 8'h30;
                    16'hC677: data_out = 8'h31;
                    16'hC678: data_out = 8'h32;
                    16'hC679: data_out = 8'h33;
                    16'hC67A: data_out = 8'h34;
                    16'hC67B: data_out = 8'h35;
                    16'hC67C: data_out = 8'h36;
                    16'hC67D: data_out = 8'h37;
                    16'hC67E: data_out = 8'h38;
                    16'hC67F: data_out = 8'h39;
                    16'hC680: data_out = 8'hC6;
                    16'hC681: data_out = 8'hC7;
                    16'hC682: data_out = 8'hC8;
                    16'hC683: data_out = 8'hC9;
                    16'hC684: data_out = 8'hCA;
                    16'hC685: data_out = 8'hCB;
                    16'hC686: data_out = 8'hCC;
                    16'hC687: data_out = 8'hCD;
                    16'hC688: data_out = 8'hCE;
                    16'hC689: data_out = 8'hCF;
                    16'hC68A: data_out = 8'hD0;
                    16'hC68B: data_out = 8'hD1;
                    16'hC68C: data_out = 8'hD2;
                    16'hC68D: data_out = 8'hD3;
                    16'hC68E: data_out = 8'hD4;
                    16'hC68F: data_out = 8'hD5;
                    16'hC690: data_out = 8'hD6;
                    16'hC691: data_out = 8'hD7;
                    16'hC692: data_out = 8'hD8;
                    16'hC693: data_out = 8'hD9;
                    16'hC694: data_out = 8'hDA;
                    16'hC695: data_out = 8'hDB;
                    16'hC696: data_out = 8'hDC;
                    16'hC697: data_out = 8'hDD;
                    16'hC698: data_out = 8'hDE;
                    16'hC699: data_out = 8'hDF;
                    16'hC69A: data_out = 8'hE0;
                    16'hC69B: data_out = 8'hE1;
                    16'hC69C: data_out = 8'hE2;
                    16'hC69D: data_out = 8'hE3;
                    16'hC69E: data_out = 8'hE4;
                    16'hC69F: data_out = 8'hE5;
                    16'hC6A0: data_out = 8'hE6;
                    16'hC6A1: data_out = 8'hE7;
                    16'hC6A2: data_out = 8'hE8;
                    16'hC6A3: data_out = 8'hE9;
                    16'hC6A4: data_out = 8'hEA;
                    16'hC6A5: data_out = 8'hEB;
                    16'hC6A6: data_out = 8'hEC;
                    16'hC6A7: data_out = 8'hED;
                    16'hC6A8: data_out = 8'hEE;
                    16'hC6A9: data_out = 8'hEF;
                    16'hC6AA: data_out = 8'hF0;
                    16'hC6AB: data_out = 8'hF1;
                    16'hC6AC: data_out = 8'hF2;
                    16'hC6AD: data_out = 8'hF3;
                    16'hC6AE: data_out = 8'hF4;
                    16'hC6AF: data_out = 8'hF5;
                    16'hC6B0: data_out = 8'hF6;
                    16'hC6B1: data_out = 8'hF7;
                    16'hC6B2: data_out = 8'hF8;
                    16'hC6B3: data_out = 8'hF9;
                    16'hC6B4: data_out = 8'hFA;
                    16'hC6B5: data_out = 8'hFB;
                    16'hC6B6: data_out = 8'hFC;
                    16'hC6B7: data_out = 8'hFD;
                    16'hC6B8: data_out = 8'hFE;
                    16'hC6B9: data_out = 8'hFF;
                    16'hC6BA: data_out = 8'h80;
                    16'hC6BB: data_out = 8'h81;
                    16'hC6BC: data_out = 8'h82;
                    16'hC6BD: data_out = 8'h83;
                    16'hC6BE: data_out = 8'h84;
                    16'hC6BF: data_out = 8'h85;
                    16'hC6C0: data_out = 8'h86;
                    16'hC6C1: data_out = 8'h87;
                    16'hC6C2: data_out = 8'h88;
                    16'hC6C3: data_out = 8'h89;
                    16'hC6C4: data_out = 8'h8A;
                    16'hC6C5: data_out = 8'h8B;
                    16'hC6C6: data_out = 8'h8C;
                    16'hC6C7: data_out = 8'h8D;
                    16'hC6C8: data_out = 8'h8E;
                    16'hC6C9: data_out = 8'h8F;
                    16'hC6CA: data_out = 8'h90;
                    16'hC6CB: data_out = 8'h91;
                    16'hC6CC: data_out = 8'h92;
                    16'hC6CD: data_out = 8'h93;
                    16'hC6CE: data_out = 8'h94;
                    16'hC6CF: data_out = 8'h95;
                    16'hC6D0: data_out = 8'h96;
                    16'hC6D1: data_out = 8'h97;
                    16'hC6D2: data_out = 8'h98;
                    16'hC6D3: data_out = 8'h99;
                    16'hC6D4: data_out = 8'h9A;
                    16'hC6D5: data_out = 8'h9B;
                    16'hC6D6: data_out = 8'h9C;
                    16'hC6D7: data_out = 8'h9D;
                    16'hC6D8: data_out = 8'h9E;
                    16'hC6D9: data_out = 8'h9F;
                    16'hC6DA: data_out = 8'hA0;
                    16'hC6DB: data_out = 8'hA1;
                    16'hC6DC: data_out = 8'hA2;
                    16'hC6DD: data_out = 8'hA3;
                    16'hC6DE: data_out = 8'hA4;
                    16'hC6DF: data_out = 8'hA5;
                    16'hC6E0: data_out = 8'hA6;
                    16'hC6E1: data_out = 8'hA7;
                    16'hC6E2: data_out = 8'hA8;
                    16'hC6E3: data_out = 8'hA9;
                    16'hC6E4: data_out = 8'hAA;
                    16'hC6E5: data_out = 8'hAB;
                    16'hC6E6: data_out = 8'hAC;
                    16'hC6E7: data_out = 8'hAD;
                    16'hC6E8: data_out = 8'hAE;
                    16'hC6E9: data_out = 8'hAF;
                    16'hC6EA: data_out = 8'hB0;
                    16'hC6EB: data_out = 8'hB1;
                    16'hC6EC: data_out = 8'hB2;
                    16'hC6ED: data_out = 8'hB3;
                    16'hC6EE: data_out = 8'hB4;
                    16'hC6EF: data_out = 8'hB5;
                    16'hC6F0: data_out = 8'hB6;
                    16'hC6F1: data_out = 8'hB7;
                    16'hC6F2: data_out = 8'hB8;
                    16'hC6F3: data_out = 8'hB9;
                    16'hC6F4: data_out = 8'hBA;
                    16'hC6F5: data_out = 8'hBB;
                    16'hC6F6: data_out = 8'hBC;
                    16'hC6F7: data_out = 8'hBD;
                    16'hC6F8: data_out = 8'hBE;
                    16'hC6F9: data_out = 8'hBF;
                    16'hC6FA: data_out = 8'hC0;
                    16'hC6FB: data_out = 8'hC1;
                    16'hC6FC: data_out = 8'hC2;
                    16'hC6FD: data_out = 8'hC3;
                    16'hC6FE: data_out = 8'hC4;
                    16'hC6FF: data_out = 8'hC5;
                    16'hC700: data_out = 8'hC7;
                    16'hC701: data_out = 8'hC6;
                    16'hC702: data_out = 8'hC5;
                    16'hC703: data_out = 8'hC4;
                    16'hC704: data_out = 8'hC3;
                    16'hC705: data_out = 8'hC2;
                    16'hC706: data_out = 8'hC1;
                    16'hC707: data_out = 8'hC0;
                    16'hC708: data_out = 8'hBF;
                    16'hC709: data_out = 8'hBE;
                    16'hC70A: data_out = 8'hBD;
                    16'hC70B: data_out = 8'hBC;
                    16'hC70C: data_out = 8'hBB;
                    16'hC70D: data_out = 8'hBA;
                    16'hC70E: data_out = 8'hB9;
                    16'hC70F: data_out = 8'hB8;
                    16'hC710: data_out = 8'hB7;
                    16'hC711: data_out = 8'hB6;
                    16'hC712: data_out = 8'hB5;
                    16'hC713: data_out = 8'hB4;
                    16'hC714: data_out = 8'hB3;
                    16'hC715: data_out = 8'hB2;
                    16'hC716: data_out = 8'hB1;
                    16'hC717: data_out = 8'hB0;
                    16'hC718: data_out = 8'hAF;
                    16'hC719: data_out = 8'hAE;
                    16'hC71A: data_out = 8'hAD;
                    16'hC71B: data_out = 8'hAC;
                    16'hC71C: data_out = 8'hAB;
                    16'hC71D: data_out = 8'hAA;
                    16'hC71E: data_out = 8'hA9;
                    16'hC71F: data_out = 8'hA8;
                    16'hC720: data_out = 8'hA7;
                    16'hC721: data_out = 8'hA6;
                    16'hC722: data_out = 8'hA5;
                    16'hC723: data_out = 8'hA4;
                    16'hC724: data_out = 8'hA3;
                    16'hC725: data_out = 8'hA2;
                    16'hC726: data_out = 8'hA1;
                    16'hC727: data_out = 8'hA0;
                    16'hC728: data_out = 8'h9F;
                    16'hC729: data_out = 8'h9E;
                    16'hC72A: data_out = 8'h9D;
                    16'hC72B: data_out = 8'h9C;
                    16'hC72C: data_out = 8'h9B;
                    16'hC72D: data_out = 8'h9A;
                    16'hC72E: data_out = 8'h99;
                    16'hC72F: data_out = 8'h98;
                    16'hC730: data_out = 8'h97;
                    16'hC731: data_out = 8'h96;
                    16'hC732: data_out = 8'h95;
                    16'hC733: data_out = 8'h94;
                    16'hC734: data_out = 8'h93;
                    16'hC735: data_out = 8'h92;
                    16'hC736: data_out = 8'h91;
                    16'hC737: data_out = 8'h90;
                    16'hC738: data_out = 8'h8F;
                    16'hC739: data_out = 8'h8E;
                    16'hC73A: data_out = 8'h8D;
                    16'hC73B: data_out = 8'h8C;
                    16'hC73C: data_out = 8'h8B;
                    16'hC73D: data_out = 8'h8A;
                    16'hC73E: data_out = 8'h89;
                    16'hC73F: data_out = 8'h88;
                    16'hC740: data_out = 8'h87;
                    16'hC741: data_out = 8'h86;
                    16'hC742: data_out = 8'h85;
                    16'hC743: data_out = 8'h84;
                    16'hC744: data_out = 8'h83;
                    16'hC745: data_out = 8'h82;
                    16'hC746: data_out = 8'h81;
                    16'hC747: data_out = 8'h0;
                    16'hC748: data_out = 8'h1;
                    16'hC749: data_out = 8'h2;
                    16'hC74A: data_out = 8'h3;
                    16'hC74B: data_out = 8'h4;
                    16'hC74C: data_out = 8'h5;
                    16'hC74D: data_out = 8'h6;
                    16'hC74E: data_out = 8'h7;
                    16'hC74F: data_out = 8'h8;
                    16'hC750: data_out = 8'h9;
                    16'hC751: data_out = 8'hA;
                    16'hC752: data_out = 8'hB;
                    16'hC753: data_out = 8'hC;
                    16'hC754: data_out = 8'hD;
                    16'hC755: data_out = 8'hE;
                    16'hC756: data_out = 8'hF;
                    16'hC757: data_out = 8'h10;
                    16'hC758: data_out = 8'h11;
                    16'hC759: data_out = 8'h12;
                    16'hC75A: data_out = 8'h13;
                    16'hC75B: data_out = 8'h14;
                    16'hC75C: data_out = 8'h15;
                    16'hC75D: data_out = 8'h16;
                    16'hC75E: data_out = 8'h17;
                    16'hC75F: data_out = 8'h18;
                    16'hC760: data_out = 8'h19;
                    16'hC761: data_out = 8'h1A;
                    16'hC762: data_out = 8'h1B;
                    16'hC763: data_out = 8'h1C;
                    16'hC764: data_out = 8'h1D;
                    16'hC765: data_out = 8'h1E;
                    16'hC766: data_out = 8'h1F;
                    16'hC767: data_out = 8'h20;
                    16'hC768: data_out = 8'h21;
                    16'hC769: data_out = 8'h22;
                    16'hC76A: data_out = 8'h23;
                    16'hC76B: data_out = 8'h24;
                    16'hC76C: data_out = 8'h25;
                    16'hC76D: data_out = 8'h26;
                    16'hC76E: data_out = 8'h27;
                    16'hC76F: data_out = 8'h28;
                    16'hC770: data_out = 8'h29;
                    16'hC771: data_out = 8'h2A;
                    16'hC772: data_out = 8'h2B;
                    16'hC773: data_out = 8'h2C;
                    16'hC774: data_out = 8'h2D;
                    16'hC775: data_out = 8'h2E;
                    16'hC776: data_out = 8'h2F;
                    16'hC777: data_out = 8'h30;
                    16'hC778: data_out = 8'h31;
                    16'hC779: data_out = 8'h32;
                    16'hC77A: data_out = 8'h33;
                    16'hC77B: data_out = 8'h34;
                    16'hC77C: data_out = 8'h35;
                    16'hC77D: data_out = 8'h36;
                    16'hC77E: data_out = 8'h37;
                    16'hC77F: data_out = 8'h38;
                    16'hC780: data_out = 8'hC7;
                    16'hC781: data_out = 8'hC8;
                    16'hC782: data_out = 8'hC9;
                    16'hC783: data_out = 8'hCA;
                    16'hC784: data_out = 8'hCB;
                    16'hC785: data_out = 8'hCC;
                    16'hC786: data_out = 8'hCD;
                    16'hC787: data_out = 8'hCE;
                    16'hC788: data_out = 8'hCF;
                    16'hC789: data_out = 8'hD0;
                    16'hC78A: data_out = 8'hD1;
                    16'hC78B: data_out = 8'hD2;
                    16'hC78C: data_out = 8'hD3;
                    16'hC78D: data_out = 8'hD4;
                    16'hC78E: data_out = 8'hD5;
                    16'hC78F: data_out = 8'hD6;
                    16'hC790: data_out = 8'hD7;
                    16'hC791: data_out = 8'hD8;
                    16'hC792: data_out = 8'hD9;
                    16'hC793: data_out = 8'hDA;
                    16'hC794: data_out = 8'hDB;
                    16'hC795: data_out = 8'hDC;
                    16'hC796: data_out = 8'hDD;
                    16'hC797: data_out = 8'hDE;
                    16'hC798: data_out = 8'hDF;
                    16'hC799: data_out = 8'hE0;
                    16'hC79A: data_out = 8'hE1;
                    16'hC79B: data_out = 8'hE2;
                    16'hC79C: data_out = 8'hE3;
                    16'hC79D: data_out = 8'hE4;
                    16'hC79E: data_out = 8'hE5;
                    16'hC79F: data_out = 8'hE6;
                    16'hC7A0: data_out = 8'hE7;
                    16'hC7A1: data_out = 8'hE8;
                    16'hC7A2: data_out = 8'hE9;
                    16'hC7A3: data_out = 8'hEA;
                    16'hC7A4: data_out = 8'hEB;
                    16'hC7A5: data_out = 8'hEC;
                    16'hC7A6: data_out = 8'hED;
                    16'hC7A7: data_out = 8'hEE;
                    16'hC7A8: data_out = 8'hEF;
                    16'hC7A9: data_out = 8'hF0;
                    16'hC7AA: data_out = 8'hF1;
                    16'hC7AB: data_out = 8'hF2;
                    16'hC7AC: data_out = 8'hF3;
                    16'hC7AD: data_out = 8'hF4;
                    16'hC7AE: data_out = 8'hF5;
                    16'hC7AF: data_out = 8'hF6;
                    16'hC7B0: data_out = 8'hF7;
                    16'hC7B1: data_out = 8'hF8;
                    16'hC7B2: data_out = 8'hF9;
                    16'hC7B3: data_out = 8'hFA;
                    16'hC7B4: data_out = 8'hFB;
                    16'hC7B5: data_out = 8'hFC;
                    16'hC7B6: data_out = 8'hFD;
                    16'hC7B7: data_out = 8'hFE;
                    16'hC7B8: data_out = 8'hFF;
                    16'hC7B9: data_out = 8'h80;
                    16'hC7BA: data_out = 8'h81;
                    16'hC7BB: data_out = 8'h82;
                    16'hC7BC: data_out = 8'h83;
                    16'hC7BD: data_out = 8'h84;
                    16'hC7BE: data_out = 8'h85;
                    16'hC7BF: data_out = 8'h86;
                    16'hC7C0: data_out = 8'h87;
                    16'hC7C1: data_out = 8'h88;
                    16'hC7C2: data_out = 8'h89;
                    16'hC7C3: data_out = 8'h8A;
                    16'hC7C4: data_out = 8'h8B;
                    16'hC7C5: data_out = 8'h8C;
                    16'hC7C6: data_out = 8'h8D;
                    16'hC7C7: data_out = 8'h8E;
                    16'hC7C8: data_out = 8'h8F;
                    16'hC7C9: data_out = 8'h90;
                    16'hC7CA: data_out = 8'h91;
                    16'hC7CB: data_out = 8'h92;
                    16'hC7CC: data_out = 8'h93;
                    16'hC7CD: data_out = 8'h94;
                    16'hC7CE: data_out = 8'h95;
                    16'hC7CF: data_out = 8'h96;
                    16'hC7D0: data_out = 8'h97;
                    16'hC7D1: data_out = 8'h98;
                    16'hC7D2: data_out = 8'h99;
                    16'hC7D3: data_out = 8'h9A;
                    16'hC7D4: data_out = 8'h9B;
                    16'hC7D5: data_out = 8'h9C;
                    16'hC7D6: data_out = 8'h9D;
                    16'hC7D7: data_out = 8'h9E;
                    16'hC7D8: data_out = 8'h9F;
                    16'hC7D9: data_out = 8'hA0;
                    16'hC7DA: data_out = 8'hA1;
                    16'hC7DB: data_out = 8'hA2;
                    16'hC7DC: data_out = 8'hA3;
                    16'hC7DD: data_out = 8'hA4;
                    16'hC7DE: data_out = 8'hA5;
                    16'hC7DF: data_out = 8'hA6;
                    16'hC7E0: data_out = 8'hA7;
                    16'hC7E1: data_out = 8'hA8;
                    16'hC7E2: data_out = 8'hA9;
                    16'hC7E3: data_out = 8'hAA;
                    16'hC7E4: data_out = 8'hAB;
                    16'hC7E5: data_out = 8'hAC;
                    16'hC7E6: data_out = 8'hAD;
                    16'hC7E7: data_out = 8'hAE;
                    16'hC7E8: data_out = 8'hAF;
                    16'hC7E9: data_out = 8'hB0;
                    16'hC7EA: data_out = 8'hB1;
                    16'hC7EB: data_out = 8'hB2;
                    16'hC7EC: data_out = 8'hB3;
                    16'hC7ED: data_out = 8'hB4;
                    16'hC7EE: data_out = 8'hB5;
                    16'hC7EF: data_out = 8'hB6;
                    16'hC7F0: data_out = 8'hB7;
                    16'hC7F1: data_out = 8'hB8;
                    16'hC7F2: data_out = 8'hB9;
                    16'hC7F3: data_out = 8'hBA;
                    16'hC7F4: data_out = 8'hBB;
                    16'hC7F5: data_out = 8'hBC;
                    16'hC7F6: data_out = 8'hBD;
                    16'hC7F7: data_out = 8'hBE;
                    16'hC7F8: data_out = 8'hBF;
                    16'hC7F9: data_out = 8'hC0;
                    16'hC7FA: data_out = 8'hC1;
                    16'hC7FB: data_out = 8'hC2;
                    16'hC7FC: data_out = 8'hC3;
                    16'hC7FD: data_out = 8'hC4;
                    16'hC7FE: data_out = 8'hC5;
                    16'hC7FF: data_out = 8'hC6;
                    16'hC800: data_out = 8'hC8;
                    16'hC801: data_out = 8'hC7;
                    16'hC802: data_out = 8'hC6;
                    16'hC803: data_out = 8'hC5;
                    16'hC804: data_out = 8'hC4;
                    16'hC805: data_out = 8'hC3;
                    16'hC806: data_out = 8'hC2;
                    16'hC807: data_out = 8'hC1;
                    16'hC808: data_out = 8'hC0;
                    16'hC809: data_out = 8'hBF;
                    16'hC80A: data_out = 8'hBE;
                    16'hC80B: data_out = 8'hBD;
                    16'hC80C: data_out = 8'hBC;
                    16'hC80D: data_out = 8'hBB;
                    16'hC80E: data_out = 8'hBA;
                    16'hC80F: data_out = 8'hB9;
                    16'hC810: data_out = 8'hB8;
                    16'hC811: data_out = 8'hB7;
                    16'hC812: data_out = 8'hB6;
                    16'hC813: data_out = 8'hB5;
                    16'hC814: data_out = 8'hB4;
                    16'hC815: data_out = 8'hB3;
                    16'hC816: data_out = 8'hB2;
                    16'hC817: data_out = 8'hB1;
                    16'hC818: data_out = 8'hB0;
                    16'hC819: data_out = 8'hAF;
                    16'hC81A: data_out = 8'hAE;
                    16'hC81B: data_out = 8'hAD;
                    16'hC81C: data_out = 8'hAC;
                    16'hC81D: data_out = 8'hAB;
                    16'hC81E: data_out = 8'hAA;
                    16'hC81F: data_out = 8'hA9;
                    16'hC820: data_out = 8'hA8;
                    16'hC821: data_out = 8'hA7;
                    16'hC822: data_out = 8'hA6;
                    16'hC823: data_out = 8'hA5;
                    16'hC824: data_out = 8'hA4;
                    16'hC825: data_out = 8'hA3;
                    16'hC826: data_out = 8'hA2;
                    16'hC827: data_out = 8'hA1;
                    16'hC828: data_out = 8'hA0;
                    16'hC829: data_out = 8'h9F;
                    16'hC82A: data_out = 8'h9E;
                    16'hC82B: data_out = 8'h9D;
                    16'hC82C: data_out = 8'h9C;
                    16'hC82D: data_out = 8'h9B;
                    16'hC82E: data_out = 8'h9A;
                    16'hC82F: data_out = 8'h99;
                    16'hC830: data_out = 8'h98;
                    16'hC831: data_out = 8'h97;
                    16'hC832: data_out = 8'h96;
                    16'hC833: data_out = 8'h95;
                    16'hC834: data_out = 8'h94;
                    16'hC835: data_out = 8'h93;
                    16'hC836: data_out = 8'h92;
                    16'hC837: data_out = 8'h91;
                    16'hC838: data_out = 8'h90;
                    16'hC839: data_out = 8'h8F;
                    16'hC83A: data_out = 8'h8E;
                    16'hC83B: data_out = 8'h8D;
                    16'hC83C: data_out = 8'h8C;
                    16'hC83D: data_out = 8'h8B;
                    16'hC83E: data_out = 8'h8A;
                    16'hC83F: data_out = 8'h89;
                    16'hC840: data_out = 8'h88;
                    16'hC841: data_out = 8'h87;
                    16'hC842: data_out = 8'h86;
                    16'hC843: data_out = 8'h85;
                    16'hC844: data_out = 8'h84;
                    16'hC845: data_out = 8'h83;
                    16'hC846: data_out = 8'h82;
                    16'hC847: data_out = 8'h81;
                    16'hC848: data_out = 8'h0;
                    16'hC849: data_out = 8'h1;
                    16'hC84A: data_out = 8'h2;
                    16'hC84B: data_out = 8'h3;
                    16'hC84C: data_out = 8'h4;
                    16'hC84D: data_out = 8'h5;
                    16'hC84E: data_out = 8'h6;
                    16'hC84F: data_out = 8'h7;
                    16'hC850: data_out = 8'h8;
                    16'hC851: data_out = 8'h9;
                    16'hC852: data_out = 8'hA;
                    16'hC853: data_out = 8'hB;
                    16'hC854: data_out = 8'hC;
                    16'hC855: data_out = 8'hD;
                    16'hC856: data_out = 8'hE;
                    16'hC857: data_out = 8'hF;
                    16'hC858: data_out = 8'h10;
                    16'hC859: data_out = 8'h11;
                    16'hC85A: data_out = 8'h12;
                    16'hC85B: data_out = 8'h13;
                    16'hC85C: data_out = 8'h14;
                    16'hC85D: data_out = 8'h15;
                    16'hC85E: data_out = 8'h16;
                    16'hC85F: data_out = 8'h17;
                    16'hC860: data_out = 8'h18;
                    16'hC861: data_out = 8'h19;
                    16'hC862: data_out = 8'h1A;
                    16'hC863: data_out = 8'h1B;
                    16'hC864: data_out = 8'h1C;
                    16'hC865: data_out = 8'h1D;
                    16'hC866: data_out = 8'h1E;
                    16'hC867: data_out = 8'h1F;
                    16'hC868: data_out = 8'h20;
                    16'hC869: data_out = 8'h21;
                    16'hC86A: data_out = 8'h22;
                    16'hC86B: data_out = 8'h23;
                    16'hC86C: data_out = 8'h24;
                    16'hC86D: data_out = 8'h25;
                    16'hC86E: data_out = 8'h26;
                    16'hC86F: data_out = 8'h27;
                    16'hC870: data_out = 8'h28;
                    16'hC871: data_out = 8'h29;
                    16'hC872: data_out = 8'h2A;
                    16'hC873: data_out = 8'h2B;
                    16'hC874: data_out = 8'h2C;
                    16'hC875: data_out = 8'h2D;
                    16'hC876: data_out = 8'h2E;
                    16'hC877: data_out = 8'h2F;
                    16'hC878: data_out = 8'h30;
                    16'hC879: data_out = 8'h31;
                    16'hC87A: data_out = 8'h32;
                    16'hC87B: data_out = 8'h33;
                    16'hC87C: data_out = 8'h34;
                    16'hC87D: data_out = 8'h35;
                    16'hC87E: data_out = 8'h36;
                    16'hC87F: data_out = 8'h37;
                    16'hC880: data_out = 8'hC8;
                    16'hC881: data_out = 8'hC9;
                    16'hC882: data_out = 8'hCA;
                    16'hC883: data_out = 8'hCB;
                    16'hC884: data_out = 8'hCC;
                    16'hC885: data_out = 8'hCD;
                    16'hC886: data_out = 8'hCE;
                    16'hC887: data_out = 8'hCF;
                    16'hC888: data_out = 8'hD0;
                    16'hC889: data_out = 8'hD1;
                    16'hC88A: data_out = 8'hD2;
                    16'hC88B: data_out = 8'hD3;
                    16'hC88C: data_out = 8'hD4;
                    16'hC88D: data_out = 8'hD5;
                    16'hC88E: data_out = 8'hD6;
                    16'hC88F: data_out = 8'hD7;
                    16'hC890: data_out = 8'hD8;
                    16'hC891: data_out = 8'hD9;
                    16'hC892: data_out = 8'hDA;
                    16'hC893: data_out = 8'hDB;
                    16'hC894: data_out = 8'hDC;
                    16'hC895: data_out = 8'hDD;
                    16'hC896: data_out = 8'hDE;
                    16'hC897: data_out = 8'hDF;
                    16'hC898: data_out = 8'hE0;
                    16'hC899: data_out = 8'hE1;
                    16'hC89A: data_out = 8'hE2;
                    16'hC89B: data_out = 8'hE3;
                    16'hC89C: data_out = 8'hE4;
                    16'hC89D: data_out = 8'hE5;
                    16'hC89E: data_out = 8'hE6;
                    16'hC89F: data_out = 8'hE7;
                    16'hC8A0: data_out = 8'hE8;
                    16'hC8A1: data_out = 8'hE9;
                    16'hC8A2: data_out = 8'hEA;
                    16'hC8A3: data_out = 8'hEB;
                    16'hC8A4: data_out = 8'hEC;
                    16'hC8A5: data_out = 8'hED;
                    16'hC8A6: data_out = 8'hEE;
                    16'hC8A7: data_out = 8'hEF;
                    16'hC8A8: data_out = 8'hF0;
                    16'hC8A9: data_out = 8'hF1;
                    16'hC8AA: data_out = 8'hF2;
                    16'hC8AB: data_out = 8'hF3;
                    16'hC8AC: data_out = 8'hF4;
                    16'hC8AD: data_out = 8'hF5;
                    16'hC8AE: data_out = 8'hF6;
                    16'hC8AF: data_out = 8'hF7;
                    16'hC8B0: data_out = 8'hF8;
                    16'hC8B1: data_out = 8'hF9;
                    16'hC8B2: data_out = 8'hFA;
                    16'hC8B3: data_out = 8'hFB;
                    16'hC8B4: data_out = 8'hFC;
                    16'hC8B5: data_out = 8'hFD;
                    16'hC8B6: data_out = 8'hFE;
                    16'hC8B7: data_out = 8'hFF;
                    16'hC8B8: data_out = 8'h80;
                    16'hC8B9: data_out = 8'h81;
                    16'hC8BA: data_out = 8'h82;
                    16'hC8BB: data_out = 8'h83;
                    16'hC8BC: data_out = 8'h84;
                    16'hC8BD: data_out = 8'h85;
                    16'hC8BE: data_out = 8'h86;
                    16'hC8BF: data_out = 8'h87;
                    16'hC8C0: data_out = 8'h88;
                    16'hC8C1: data_out = 8'h89;
                    16'hC8C2: data_out = 8'h8A;
                    16'hC8C3: data_out = 8'h8B;
                    16'hC8C4: data_out = 8'h8C;
                    16'hC8C5: data_out = 8'h8D;
                    16'hC8C6: data_out = 8'h8E;
                    16'hC8C7: data_out = 8'h8F;
                    16'hC8C8: data_out = 8'h90;
                    16'hC8C9: data_out = 8'h91;
                    16'hC8CA: data_out = 8'h92;
                    16'hC8CB: data_out = 8'h93;
                    16'hC8CC: data_out = 8'h94;
                    16'hC8CD: data_out = 8'h95;
                    16'hC8CE: data_out = 8'h96;
                    16'hC8CF: data_out = 8'h97;
                    16'hC8D0: data_out = 8'h98;
                    16'hC8D1: data_out = 8'h99;
                    16'hC8D2: data_out = 8'h9A;
                    16'hC8D3: data_out = 8'h9B;
                    16'hC8D4: data_out = 8'h9C;
                    16'hC8D5: data_out = 8'h9D;
                    16'hC8D6: data_out = 8'h9E;
                    16'hC8D7: data_out = 8'h9F;
                    16'hC8D8: data_out = 8'hA0;
                    16'hC8D9: data_out = 8'hA1;
                    16'hC8DA: data_out = 8'hA2;
                    16'hC8DB: data_out = 8'hA3;
                    16'hC8DC: data_out = 8'hA4;
                    16'hC8DD: data_out = 8'hA5;
                    16'hC8DE: data_out = 8'hA6;
                    16'hC8DF: data_out = 8'hA7;
                    16'hC8E0: data_out = 8'hA8;
                    16'hC8E1: data_out = 8'hA9;
                    16'hC8E2: data_out = 8'hAA;
                    16'hC8E3: data_out = 8'hAB;
                    16'hC8E4: data_out = 8'hAC;
                    16'hC8E5: data_out = 8'hAD;
                    16'hC8E6: data_out = 8'hAE;
                    16'hC8E7: data_out = 8'hAF;
                    16'hC8E8: data_out = 8'hB0;
                    16'hC8E9: data_out = 8'hB1;
                    16'hC8EA: data_out = 8'hB2;
                    16'hC8EB: data_out = 8'hB3;
                    16'hC8EC: data_out = 8'hB4;
                    16'hC8ED: data_out = 8'hB5;
                    16'hC8EE: data_out = 8'hB6;
                    16'hC8EF: data_out = 8'hB7;
                    16'hC8F0: data_out = 8'hB8;
                    16'hC8F1: data_out = 8'hB9;
                    16'hC8F2: data_out = 8'hBA;
                    16'hC8F3: data_out = 8'hBB;
                    16'hC8F4: data_out = 8'hBC;
                    16'hC8F5: data_out = 8'hBD;
                    16'hC8F6: data_out = 8'hBE;
                    16'hC8F7: data_out = 8'hBF;
                    16'hC8F8: data_out = 8'hC0;
                    16'hC8F9: data_out = 8'hC1;
                    16'hC8FA: data_out = 8'hC2;
                    16'hC8FB: data_out = 8'hC3;
                    16'hC8FC: data_out = 8'hC4;
                    16'hC8FD: data_out = 8'hC5;
                    16'hC8FE: data_out = 8'hC6;
                    16'hC8FF: data_out = 8'hC7;
                    16'hC900: data_out = 8'hC9;
                    16'hC901: data_out = 8'hC8;
                    16'hC902: data_out = 8'hC7;
                    16'hC903: data_out = 8'hC6;
                    16'hC904: data_out = 8'hC5;
                    16'hC905: data_out = 8'hC4;
                    16'hC906: data_out = 8'hC3;
                    16'hC907: data_out = 8'hC2;
                    16'hC908: data_out = 8'hC1;
                    16'hC909: data_out = 8'hC0;
                    16'hC90A: data_out = 8'hBF;
                    16'hC90B: data_out = 8'hBE;
                    16'hC90C: data_out = 8'hBD;
                    16'hC90D: data_out = 8'hBC;
                    16'hC90E: data_out = 8'hBB;
                    16'hC90F: data_out = 8'hBA;
                    16'hC910: data_out = 8'hB9;
                    16'hC911: data_out = 8'hB8;
                    16'hC912: data_out = 8'hB7;
                    16'hC913: data_out = 8'hB6;
                    16'hC914: data_out = 8'hB5;
                    16'hC915: data_out = 8'hB4;
                    16'hC916: data_out = 8'hB3;
                    16'hC917: data_out = 8'hB2;
                    16'hC918: data_out = 8'hB1;
                    16'hC919: data_out = 8'hB0;
                    16'hC91A: data_out = 8'hAF;
                    16'hC91B: data_out = 8'hAE;
                    16'hC91C: data_out = 8'hAD;
                    16'hC91D: data_out = 8'hAC;
                    16'hC91E: data_out = 8'hAB;
                    16'hC91F: data_out = 8'hAA;
                    16'hC920: data_out = 8'hA9;
                    16'hC921: data_out = 8'hA8;
                    16'hC922: data_out = 8'hA7;
                    16'hC923: data_out = 8'hA6;
                    16'hC924: data_out = 8'hA5;
                    16'hC925: data_out = 8'hA4;
                    16'hC926: data_out = 8'hA3;
                    16'hC927: data_out = 8'hA2;
                    16'hC928: data_out = 8'hA1;
                    16'hC929: data_out = 8'hA0;
                    16'hC92A: data_out = 8'h9F;
                    16'hC92B: data_out = 8'h9E;
                    16'hC92C: data_out = 8'h9D;
                    16'hC92D: data_out = 8'h9C;
                    16'hC92E: data_out = 8'h9B;
                    16'hC92F: data_out = 8'h9A;
                    16'hC930: data_out = 8'h99;
                    16'hC931: data_out = 8'h98;
                    16'hC932: data_out = 8'h97;
                    16'hC933: data_out = 8'h96;
                    16'hC934: data_out = 8'h95;
                    16'hC935: data_out = 8'h94;
                    16'hC936: data_out = 8'h93;
                    16'hC937: data_out = 8'h92;
                    16'hC938: data_out = 8'h91;
                    16'hC939: data_out = 8'h90;
                    16'hC93A: data_out = 8'h8F;
                    16'hC93B: data_out = 8'h8E;
                    16'hC93C: data_out = 8'h8D;
                    16'hC93D: data_out = 8'h8C;
                    16'hC93E: data_out = 8'h8B;
                    16'hC93F: data_out = 8'h8A;
                    16'hC940: data_out = 8'h89;
                    16'hC941: data_out = 8'h88;
                    16'hC942: data_out = 8'h87;
                    16'hC943: data_out = 8'h86;
                    16'hC944: data_out = 8'h85;
                    16'hC945: data_out = 8'h84;
                    16'hC946: data_out = 8'h83;
                    16'hC947: data_out = 8'h82;
                    16'hC948: data_out = 8'h81;
                    16'hC949: data_out = 8'h0;
                    16'hC94A: data_out = 8'h1;
                    16'hC94B: data_out = 8'h2;
                    16'hC94C: data_out = 8'h3;
                    16'hC94D: data_out = 8'h4;
                    16'hC94E: data_out = 8'h5;
                    16'hC94F: data_out = 8'h6;
                    16'hC950: data_out = 8'h7;
                    16'hC951: data_out = 8'h8;
                    16'hC952: data_out = 8'h9;
                    16'hC953: data_out = 8'hA;
                    16'hC954: data_out = 8'hB;
                    16'hC955: data_out = 8'hC;
                    16'hC956: data_out = 8'hD;
                    16'hC957: data_out = 8'hE;
                    16'hC958: data_out = 8'hF;
                    16'hC959: data_out = 8'h10;
                    16'hC95A: data_out = 8'h11;
                    16'hC95B: data_out = 8'h12;
                    16'hC95C: data_out = 8'h13;
                    16'hC95D: data_out = 8'h14;
                    16'hC95E: data_out = 8'h15;
                    16'hC95F: data_out = 8'h16;
                    16'hC960: data_out = 8'h17;
                    16'hC961: data_out = 8'h18;
                    16'hC962: data_out = 8'h19;
                    16'hC963: data_out = 8'h1A;
                    16'hC964: data_out = 8'h1B;
                    16'hC965: data_out = 8'h1C;
                    16'hC966: data_out = 8'h1D;
                    16'hC967: data_out = 8'h1E;
                    16'hC968: data_out = 8'h1F;
                    16'hC969: data_out = 8'h20;
                    16'hC96A: data_out = 8'h21;
                    16'hC96B: data_out = 8'h22;
                    16'hC96C: data_out = 8'h23;
                    16'hC96D: data_out = 8'h24;
                    16'hC96E: data_out = 8'h25;
                    16'hC96F: data_out = 8'h26;
                    16'hC970: data_out = 8'h27;
                    16'hC971: data_out = 8'h28;
                    16'hC972: data_out = 8'h29;
                    16'hC973: data_out = 8'h2A;
                    16'hC974: data_out = 8'h2B;
                    16'hC975: data_out = 8'h2C;
                    16'hC976: data_out = 8'h2D;
                    16'hC977: data_out = 8'h2E;
                    16'hC978: data_out = 8'h2F;
                    16'hC979: data_out = 8'h30;
                    16'hC97A: data_out = 8'h31;
                    16'hC97B: data_out = 8'h32;
                    16'hC97C: data_out = 8'h33;
                    16'hC97D: data_out = 8'h34;
                    16'hC97E: data_out = 8'h35;
                    16'hC97F: data_out = 8'h36;
                    16'hC980: data_out = 8'hC9;
                    16'hC981: data_out = 8'hCA;
                    16'hC982: data_out = 8'hCB;
                    16'hC983: data_out = 8'hCC;
                    16'hC984: data_out = 8'hCD;
                    16'hC985: data_out = 8'hCE;
                    16'hC986: data_out = 8'hCF;
                    16'hC987: data_out = 8'hD0;
                    16'hC988: data_out = 8'hD1;
                    16'hC989: data_out = 8'hD2;
                    16'hC98A: data_out = 8'hD3;
                    16'hC98B: data_out = 8'hD4;
                    16'hC98C: data_out = 8'hD5;
                    16'hC98D: data_out = 8'hD6;
                    16'hC98E: data_out = 8'hD7;
                    16'hC98F: data_out = 8'hD8;
                    16'hC990: data_out = 8'hD9;
                    16'hC991: data_out = 8'hDA;
                    16'hC992: data_out = 8'hDB;
                    16'hC993: data_out = 8'hDC;
                    16'hC994: data_out = 8'hDD;
                    16'hC995: data_out = 8'hDE;
                    16'hC996: data_out = 8'hDF;
                    16'hC997: data_out = 8'hE0;
                    16'hC998: data_out = 8'hE1;
                    16'hC999: data_out = 8'hE2;
                    16'hC99A: data_out = 8'hE3;
                    16'hC99B: data_out = 8'hE4;
                    16'hC99C: data_out = 8'hE5;
                    16'hC99D: data_out = 8'hE6;
                    16'hC99E: data_out = 8'hE7;
                    16'hC99F: data_out = 8'hE8;
                    16'hC9A0: data_out = 8'hE9;
                    16'hC9A1: data_out = 8'hEA;
                    16'hC9A2: data_out = 8'hEB;
                    16'hC9A3: data_out = 8'hEC;
                    16'hC9A4: data_out = 8'hED;
                    16'hC9A5: data_out = 8'hEE;
                    16'hC9A6: data_out = 8'hEF;
                    16'hC9A7: data_out = 8'hF0;
                    16'hC9A8: data_out = 8'hF1;
                    16'hC9A9: data_out = 8'hF2;
                    16'hC9AA: data_out = 8'hF3;
                    16'hC9AB: data_out = 8'hF4;
                    16'hC9AC: data_out = 8'hF5;
                    16'hC9AD: data_out = 8'hF6;
                    16'hC9AE: data_out = 8'hF7;
                    16'hC9AF: data_out = 8'hF8;
                    16'hC9B0: data_out = 8'hF9;
                    16'hC9B1: data_out = 8'hFA;
                    16'hC9B2: data_out = 8'hFB;
                    16'hC9B3: data_out = 8'hFC;
                    16'hC9B4: data_out = 8'hFD;
                    16'hC9B5: data_out = 8'hFE;
                    16'hC9B6: data_out = 8'hFF;
                    16'hC9B7: data_out = 8'h80;
                    16'hC9B8: data_out = 8'h81;
                    16'hC9B9: data_out = 8'h82;
                    16'hC9BA: data_out = 8'h83;
                    16'hC9BB: data_out = 8'h84;
                    16'hC9BC: data_out = 8'h85;
                    16'hC9BD: data_out = 8'h86;
                    16'hC9BE: data_out = 8'h87;
                    16'hC9BF: data_out = 8'h88;
                    16'hC9C0: data_out = 8'h89;
                    16'hC9C1: data_out = 8'h8A;
                    16'hC9C2: data_out = 8'h8B;
                    16'hC9C3: data_out = 8'h8C;
                    16'hC9C4: data_out = 8'h8D;
                    16'hC9C5: data_out = 8'h8E;
                    16'hC9C6: data_out = 8'h8F;
                    16'hC9C7: data_out = 8'h90;
                    16'hC9C8: data_out = 8'h91;
                    16'hC9C9: data_out = 8'h92;
                    16'hC9CA: data_out = 8'h93;
                    16'hC9CB: data_out = 8'h94;
                    16'hC9CC: data_out = 8'h95;
                    16'hC9CD: data_out = 8'h96;
                    16'hC9CE: data_out = 8'h97;
                    16'hC9CF: data_out = 8'h98;
                    16'hC9D0: data_out = 8'h99;
                    16'hC9D1: data_out = 8'h9A;
                    16'hC9D2: data_out = 8'h9B;
                    16'hC9D3: data_out = 8'h9C;
                    16'hC9D4: data_out = 8'h9D;
                    16'hC9D5: data_out = 8'h9E;
                    16'hC9D6: data_out = 8'h9F;
                    16'hC9D7: data_out = 8'hA0;
                    16'hC9D8: data_out = 8'hA1;
                    16'hC9D9: data_out = 8'hA2;
                    16'hC9DA: data_out = 8'hA3;
                    16'hC9DB: data_out = 8'hA4;
                    16'hC9DC: data_out = 8'hA5;
                    16'hC9DD: data_out = 8'hA6;
                    16'hC9DE: data_out = 8'hA7;
                    16'hC9DF: data_out = 8'hA8;
                    16'hC9E0: data_out = 8'hA9;
                    16'hC9E1: data_out = 8'hAA;
                    16'hC9E2: data_out = 8'hAB;
                    16'hC9E3: data_out = 8'hAC;
                    16'hC9E4: data_out = 8'hAD;
                    16'hC9E5: data_out = 8'hAE;
                    16'hC9E6: data_out = 8'hAF;
                    16'hC9E7: data_out = 8'hB0;
                    16'hC9E8: data_out = 8'hB1;
                    16'hC9E9: data_out = 8'hB2;
                    16'hC9EA: data_out = 8'hB3;
                    16'hC9EB: data_out = 8'hB4;
                    16'hC9EC: data_out = 8'hB5;
                    16'hC9ED: data_out = 8'hB6;
                    16'hC9EE: data_out = 8'hB7;
                    16'hC9EF: data_out = 8'hB8;
                    16'hC9F0: data_out = 8'hB9;
                    16'hC9F1: data_out = 8'hBA;
                    16'hC9F2: data_out = 8'hBB;
                    16'hC9F3: data_out = 8'hBC;
                    16'hC9F4: data_out = 8'hBD;
                    16'hC9F5: data_out = 8'hBE;
                    16'hC9F6: data_out = 8'hBF;
                    16'hC9F7: data_out = 8'hC0;
                    16'hC9F8: data_out = 8'hC1;
                    16'hC9F9: data_out = 8'hC2;
                    16'hC9FA: data_out = 8'hC3;
                    16'hC9FB: data_out = 8'hC4;
                    16'hC9FC: data_out = 8'hC5;
                    16'hC9FD: data_out = 8'hC6;
                    16'hC9FE: data_out = 8'hC7;
                    16'hC9FF: data_out = 8'hC8;
                    16'hCA00: data_out = 8'hCA;
                    16'hCA01: data_out = 8'hC9;
                    16'hCA02: data_out = 8'hC8;
                    16'hCA03: data_out = 8'hC7;
                    16'hCA04: data_out = 8'hC6;
                    16'hCA05: data_out = 8'hC5;
                    16'hCA06: data_out = 8'hC4;
                    16'hCA07: data_out = 8'hC3;
                    16'hCA08: data_out = 8'hC2;
                    16'hCA09: data_out = 8'hC1;
                    16'hCA0A: data_out = 8'hC0;
                    16'hCA0B: data_out = 8'hBF;
                    16'hCA0C: data_out = 8'hBE;
                    16'hCA0D: data_out = 8'hBD;
                    16'hCA0E: data_out = 8'hBC;
                    16'hCA0F: data_out = 8'hBB;
                    16'hCA10: data_out = 8'hBA;
                    16'hCA11: data_out = 8'hB9;
                    16'hCA12: data_out = 8'hB8;
                    16'hCA13: data_out = 8'hB7;
                    16'hCA14: data_out = 8'hB6;
                    16'hCA15: data_out = 8'hB5;
                    16'hCA16: data_out = 8'hB4;
                    16'hCA17: data_out = 8'hB3;
                    16'hCA18: data_out = 8'hB2;
                    16'hCA19: data_out = 8'hB1;
                    16'hCA1A: data_out = 8'hB0;
                    16'hCA1B: data_out = 8'hAF;
                    16'hCA1C: data_out = 8'hAE;
                    16'hCA1D: data_out = 8'hAD;
                    16'hCA1E: data_out = 8'hAC;
                    16'hCA1F: data_out = 8'hAB;
                    16'hCA20: data_out = 8'hAA;
                    16'hCA21: data_out = 8'hA9;
                    16'hCA22: data_out = 8'hA8;
                    16'hCA23: data_out = 8'hA7;
                    16'hCA24: data_out = 8'hA6;
                    16'hCA25: data_out = 8'hA5;
                    16'hCA26: data_out = 8'hA4;
                    16'hCA27: data_out = 8'hA3;
                    16'hCA28: data_out = 8'hA2;
                    16'hCA29: data_out = 8'hA1;
                    16'hCA2A: data_out = 8'hA0;
                    16'hCA2B: data_out = 8'h9F;
                    16'hCA2C: data_out = 8'h9E;
                    16'hCA2D: data_out = 8'h9D;
                    16'hCA2E: data_out = 8'h9C;
                    16'hCA2F: data_out = 8'h9B;
                    16'hCA30: data_out = 8'h9A;
                    16'hCA31: data_out = 8'h99;
                    16'hCA32: data_out = 8'h98;
                    16'hCA33: data_out = 8'h97;
                    16'hCA34: data_out = 8'h96;
                    16'hCA35: data_out = 8'h95;
                    16'hCA36: data_out = 8'h94;
                    16'hCA37: data_out = 8'h93;
                    16'hCA38: data_out = 8'h92;
                    16'hCA39: data_out = 8'h91;
                    16'hCA3A: data_out = 8'h90;
                    16'hCA3B: data_out = 8'h8F;
                    16'hCA3C: data_out = 8'h8E;
                    16'hCA3D: data_out = 8'h8D;
                    16'hCA3E: data_out = 8'h8C;
                    16'hCA3F: data_out = 8'h8B;
                    16'hCA40: data_out = 8'h8A;
                    16'hCA41: data_out = 8'h89;
                    16'hCA42: data_out = 8'h88;
                    16'hCA43: data_out = 8'h87;
                    16'hCA44: data_out = 8'h86;
                    16'hCA45: data_out = 8'h85;
                    16'hCA46: data_out = 8'h84;
                    16'hCA47: data_out = 8'h83;
                    16'hCA48: data_out = 8'h82;
                    16'hCA49: data_out = 8'h81;
                    16'hCA4A: data_out = 8'h0;
                    16'hCA4B: data_out = 8'h1;
                    16'hCA4C: data_out = 8'h2;
                    16'hCA4D: data_out = 8'h3;
                    16'hCA4E: data_out = 8'h4;
                    16'hCA4F: data_out = 8'h5;
                    16'hCA50: data_out = 8'h6;
                    16'hCA51: data_out = 8'h7;
                    16'hCA52: data_out = 8'h8;
                    16'hCA53: data_out = 8'h9;
                    16'hCA54: data_out = 8'hA;
                    16'hCA55: data_out = 8'hB;
                    16'hCA56: data_out = 8'hC;
                    16'hCA57: data_out = 8'hD;
                    16'hCA58: data_out = 8'hE;
                    16'hCA59: data_out = 8'hF;
                    16'hCA5A: data_out = 8'h10;
                    16'hCA5B: data_out = 8'h11;
                    16'hCA5C: data_out = 8'h12;
                    16'hCA5D: data_out = 8'h13;
                    16'hCA5E: data_out = 8'h14;
                    16'hCA5F: data_out = 8'h15;
                    16'hCA60: data_out = 8'h16;
                    16'hCA61: data_out = 8'h17;
                    16'hCA62: data_out = 8'h18;
                    16'hCA63: data_out = 8'h19;
                    16'hCA64: data_out = 8'h1A;
                    16'hCA65: data_out = 8'h1B;
                    16'hCA66: data_out = 8'h1C;
                    16'hCA67: data_out = 8'h1D;
                    16'hCA68: data_out = 8'h1E;
                    16'hCA69: data_out = 8'h1F;
                    16'hCA6A: data_out = 8'h20;
                    16'hCA6B: data_out = 8'h21;
                    16'hCA6C: data_out = 8'h22;
                    16'hCA6D: data_out = 8'h23;
                    16'hCA6E: data_out = 8'h24;
                    16'hCA6F: data_out = 8'h25;
                    16'hCA70: data_out = 8'h26;
                    16'hCA71: data_out = 8'h27;
                    16'hCA72: data_out = 8'h28;
                    16'hCA73: data_out = 8'h29;
                    16'hCA74: data_out = 8'h2A;
                    16'hCA75: data_out = 8'h2B;
                    16'hCA76: data_out = 8'h2C;
                    16'hCA77: data_out = 8'h2D;
                    16'hCA78: data_out = 8'h2E;
                    16'hCA79: data_out = 8'h2F;
                    16'hCA7A: data_out = 8'h30;
                    16'hCA7B: data_out = 8'h31;
                    16'hCA7C: data_out = 8'h32;
                    16'hCA7D: data_out = 8'h33;
                    16'hCA7E: data_out = 8'h34;
                    16'hCA7F: data_out = 8'h35;
                    16'hCA80: data_out = 8'hCA;
                    16'hCA81: data_out = 8'hCB;
                    16'hCA82: data_out = 8'hCC;
                    16'hCA83: data_out = 8'hCD;
                    16'hCA84: data_out = 8'hCE;
                    16'hCA85: data_out = 8'hCF;
                    16'hCA86: data_out = 8'hD0;
                    16'hCA87: data_out = 8'hD1;
                    16'hCA88: data_out = 8'hD2;
                    16'hCA89: data_out = 8'hD3;
                    16'hCA8A: data_out = 8'hD4;
                    16'hCA8B: data_out = 8'hD5;
                    16'hCA8C: data_out = 8'hD6;
                    16'hCA8D: data_out = 8'hD7;
                    16'hCA8E: data_out = 8'hD8;
                    16'hCA8F: data_out = 8'hD9;
                    16'hCA90: data_out = 8'hDA;
                    16'hCA91: data_out = 8'hDB;
                    16'hCA92: data_out = 8'hDC;
                    16'hCA93: data_out = 8'hDD;
                    16'hCA94: data_out = 8'hDE;
                    16'hCA95: data_out = 8'hDF;
                    16'hCA96: data_out = 8'hE0;
                    16'hCA97: data_out = 8'hE1;
                    16'hCA98: data_out = 8'hE2;
                    16'hCA99: data_out = 8'hE3;
                    16'hCA9A: data_out = 8'hE4;
                    16'hCA9B: data_out = 8'hE5;
                    16'hCA9C: data_out = 8'hE6;
                    16'hCA9D: data_out = 8'hE7;
                    16'hCA9E: data_out = 8'hE8;
                    16'hCA9F: data_out = 8'hE9;
                    16'hCAA0: data_out = 8'hEA;
                    16'hCAA1: data_out = 8'hEB;
                    16'hCAA2: data_out = 8'hEC;
                    16'hCAA3: data_out = 8'hED;
                    16'hCAA4: data_out = 8'hEE;
                    16'hCAA5: data_out = 8'hEF;
                    16'hCAA6: data_out = 8'hF0;
                    16'hCAA7: data_out = 8'hF1;
                    16'hCAA8: data_out = 8'hF2;
                    16'hCAA9: data_out = 8'hF3;
                    16'hCAAA: data_out = 8'hF4;
                    16'hCAAB: data_out = 8'hF5;
                    16'hCAAC: data_out = 8'hF6;
                    16'hCAAD: data_out = 8'hF7;
                    16'hCAAE: data_out = 8'hF8;
                    16'hCAAF: data_out = 8'hF9;
                    16'hCAB0: data_out = 8'hFA;
                    16'hCAB1: data_out = 8'hFB;
                    16'hCAB2: data_out = 8'hFC;
                    16'hCAB3: data_out = 8'hFD;
                    16'hCAB4: data_out = 8'hFE;
                    16'hCAB5: data_out = 8'hFF;
                    16'hCAB6: data_out = 8'h80;
                    16'hCAB7: data_out = 8'h81;
                    16'hCAB8: data_out = 8'h82;
                    16'hCAB9: data_out = 8'h83;
                    16'hCABA: data_out = 8'h84;
                    16'hCABB: data_out = 8'h85;
                    16'hCABC: data_out = 8'h86;
                    16'hCABD: data_out = 8'h87;
                    16'hCABE: data_out = 8'h88;
                    16'hCABF: data_out = 8'h89;
                    16'hCAC0: data_out = 8'h8A;
                    16'hCAC1: data_out = 8'h8B;
                    16'hCAC2: data_out = 8'h8C;
                    16'hCAC3: data_out = 8'h8D;
                    16'hCAC4: data_out = 8'h8E;
                    16'hCAC5: data_out = 8'h8F;
                    16'hCAC6: data_out = 8'h90;
                    16'hCAC7: data_out = 8'h91;
                    16'hCAC8: data_out = 8'h92;
                    16'hCAC9: data_out = 8'h93;
                    16'hCACA: data_out = 8'h94;
                    16'hCACB: data_out = 8'h95;
                    16'hCACC: data_out = 8'h96;
                    16'hCACD: data_out = 8'h97;
                    16'hCACE: data_out = 8'h98;
                    16'hCACF: data_out = 8'h99;
                    16'hCAD0: data_out = 8'h9A;
                    16'hCAD1: data_out = 8'h9B;
                    16'hCAD2: data_out = 8'h9C;
                    16'hCAD3: data_out = 8'h9D;
                    16'hCAD4: data_out = 8'h9E;
                    16'hCAD5: data_out = 8'h9F;
                    16'hCAD6: data_out = 8'hA0;
                    16'hCAD7: data_out = 8'hA1;
                    16'hCAD8: data_out = 8'hA2;
                    16'hCAD9: data_out = 8'hA3;
                    16'hCADA: data_out = 8'hA4;
                    16'hCADB: data_out = 8'hA5;
                    16'hCADC: data_out = 8'hA6;
                    16'hCADD: data_out = 8'hA7;
                    16'hCADE: data_out = 8'hA8;
                    16'hCADF: data_out = 8'hA9;
                    16'hCAE0: data_out = 8'hAA;
                    16'hCAE1: data_out = 8'hAB;
                    16'hCAE2: data_out = 8'hAC;
                    16'hCAE3: data_out = 8'hAD;
                    16'hCAE4: data_out = 8'hAE;
                    16'hCAE5: data_out = 8'hAF;
                    16'hCAE6: data_out = 8'hB0;
                    16'hCAE7: data_out = 8'hB1;
                    16'hCAE8: data_out = 8'hB2;
                    16'hCAE9: data_out = 8'hB3;
                    16'hCAEA: data_out = 8'hB4;
                    16'hCAEB: data_out = 8'hB5;
                    16'hCAEC: data_out = 8'hB6;
                    16'hCAED: data_out = 8'hB7;
                    16'hCAEE: data_out = 8'hB8;
                    16'hCAEF: data_out = 8'hB9;
                    16'hCAF0: data_out = 8'hBA;
                    16'hCAF1: data_out = 8'hBB;
                    16'hCAF2: data_out = 8'hBC;
                    16'hCAF3: data_out = 8'hBD;
                    16'hCAF4: data_out = 8'hBE;
                    16'hCAF5: data_out = 8'hBF;
                    16'hCAF6: data_out = 8'hC0;
                    16'hCAF7: data_out = 8'hC1;
                    16'hCAF8: data_out = 8'hC2;
                    16'hCAF9: data_out = 8'hC3;
                    16'hCAFA: data_out = 8'hC4;
                    16'hCAFB: data_out = 8'hC5;
                    16'hCAFC: data_out = 8'hC6;
                    16'hCAFD: data_out = 8'hC7;
                    16'hCAFE: data_out = 8'hC8;
                    16'hCAFF: data_out = 8'hC9;
                    16'hCB00: data_out = 8'hCB;
                    16'hCB01: data_out = 8'hCA;
                    16'hCB02: data_out = 8'hC9;
                    16'hCB03: data_out = 8'hC8;
                    16'hCB04: data_out = 8'hC7;
                    16'hCB05: data_out = 8'hC6;
                    16'hCB06: data_out = 8'hC5;
                    16'hCB07: data_out = 8'hC4;
                    16'hCB08: data_out = 8'hC3;
                    16'hCB09: data_out = 8'hC2;
                    16'hCB0A: data_out = 8'hC1;
                    16'hCB0B: data_out = 8'hC0;
                    16'hCB0C: data_out = 8'hBF;
                    16'hCB0D: data_out = 8'hBE;
                    16'hCB0E: data_out = 8'hBD;
                    16'hCB0F: data_out = 8'hBC;
                    16'hCB10: data_out = 8'hBB;
                    16'hCB11: data_out = 8'hBA;
                    16'hCB12: data_out = 8'hB9;
                    16'hCB13: data_out = 8'hB8;
                    16'hCB14: data_out = 8'hB7;
                    16'hCB15: data_out = 8'hB6;
                    16'hCB16: data_out = 8'hB5;
                    16'hCB17: data_out = 8'hB4;
                    16'hCB18: data_out = 8'hB3;
                    16'hCB19: data_out = 8'hB2;
                    16'hCB1A: data_out = 8'hB1;
                    16'hCB1B: data_out = 8'hB0;
                    16'hCB1C: data_out = 8'hAF;
                    16'hCB1D: data_out = 8'hAE;
                    16'hCB1E: data_out = 8'hAD;
                    16'hCB1F: data_out = 8'hAC;
                    16'hCB20: data_out = 8'hAB;
                    16'hCB21: data_out = 8'hAA;
                    16'hCB22: data_out = 8'hA9;
                    16'hCB23: data_out = 8'hA8;
                    16'hCB24: data_out = 8'hA7;
                    16'hCB25: data_out = 8'hA6;
                    16'hCB26: data_out = 8'hA5;
                    16'hCB27: data_out = 8'hA4;
                    16'hCB28: data_out = 8'hA3;
                    16'hCB29: data_out = 8'hA2;
                    16'hCB2A: data_out = 8'hA1;
                    16'hCB2B: data_out = 8'hA0;
                    16'hCB2C: data_out = 8'h9F;
                    16'hCB2D: data_out = 8'h9E;
                    16'hCB2E: data_out = 8'h9D;
                    16'hCB2F: data_out = 8'h9C;
                    16'hCB30: data_out = 8'h9B;
                    16'hCB31: data_out = 8'h9A;
                    16'hCB32: data_out = 8'h99;
                    16'hCB33: data_out = 8'h98;
                    16'hCB34: data_out = 8'h97;
                    16'hCB35: data_out = 8'h96;
                    16'hCB36: data_out = 8'h95;
                    16'hCB37: data_out = 8'h94;
                    16'hCB38: data_out = 8'h93;
                    16'hCB39: data_out = 8'h92;
                    16'hCB3A: data_out = 8'h91;
                    16'hCB3B: data_out = 8'h90;
                    16'hCB3C: data_out = 8'h8F;
                    16'hCB3D: data_out = 8'h8E;
                    16'hCB3E: data_out = 8'h8D;
                    16'hCB3F: data_out = 8'h8C;
                    16'hCB40: data_out = 8'h8B;
                    16'hCB41: data_out = 8'h8A;
                    16'hCB42: data_out = 8'h89;
                    16'hCB43: data_out = 8'h88;
                    16'hCB44: data_out = 8'h87;
                    16'hCB45: data_out = 8'h86;
                    16'hCB46: data_out = 8'h85;
                    16'hCB47: data_out = 8'h84;
                    16'hCB48: data_out = 8'h83;
                    16'hCB49: data_out = 8'h82;
                    16'hCB4A: data_out = 8'h81;
                    16'hCB4B: data_out = 8'h0;
                    16'hCB4C: data_out = 8'h1;
                    16'hCB4D: data_out = 8'h2;
                    16'hCB4E: data_out = 8'h3;
                    16'hCB4F: data_out = 8'h4;
                    16'hCB50: data_out = 8'h5;
                    16'hCB51: data_out = 8'h6;
                    16'hCB52: data_out = 8'h7;
                    16'hCB53: data_out = 8'h8;
                    16'hCB54: data_out = 8'h9;
                    16'hCB55: data_out = 8'hA;
                    16'hCB56: data_out = 8'hB;
                    16'hCB57: data_out = 8'hC;
                    16'hCB58: data_out = 8'hD;
                    16'hCB59: data_out = 8'hE;
                    16'hCB5A: data_out = 8'hF;
                    16'hCB5B: data_out = 8'h10;
                    16'hCB5C: data_out = 8'h11;
                    16'hCB5D: data_out = 8'h12;
                    16'hCB5E: data_out = 8'h13;
                    16'hCB5F: data_out = 8'h14;
                    16'hCB60: data_out = 8'h15;
                    16'hCB61: data_out = 8'h16;
                    16'hCB62: data_out = 8'h17;
                    16'hCB63: data_out = 8'h18;
                    16'hCB64: data_out = 8'h19;
                    16'hCB65: data_out = 8'h1A;
                    16'hCB66: data_out = 8'h1B;
                    16'hCB67: data_out = 8'h1C;
                    16'hCB68: data_out = 8'h1D;
                    16'hCB69: data_out = 8'h1E;
                    16'hCB6A: data_out = 8'h1F;
                    16'hCB6B: data_out = 8'h20;
                    16'hCB6C: data_out = 8'h21;
                    16'hCB6D: data_out = 8'h22;
                    16'hCB6E: data_out = 8'h23;
                    16'hCB6F: data_out = 8'h24;
                    16'hCB70: data_out = 8'h25;
                    16'hCB71: data_out = 8'h26;
                    16'hCB72: data_out = 8'h27;
                    16'hCB73: data_out = 8'h28;
                    16'hCB74: data_out = 8'h29;
                    16'hCB75: data_out = 8'h2A;
                    16'hCB76: data_out = 8'h2B;
                    16'hCB77: data_out = 8'h2C;
                    16'hCB78: data_out = 8'h2D;
                    16'hCB79: data_out = 8'h2E;
                    16'hCB7A: data_out = 8'h2F;
                    16'hCB7B: data_out = 8'h30;
                    16'hCB7C: data_out = 8'h31;
                    16'hCB7D: data_out = 8'h32;
                    16'hCB7E: data_out = 8'h33;
                    16'hCB7F: data_out = 8'h34;
                    16'hCB80: data_out = 8'hCB;
                    16'hCB81: data_out = 8'hCC;
                    16'hCB82: data_out = 8'hCD;
                    16'hCB83: data_out = 8'hCE;
                    16'hCB84: data_out = 8'hCF;
                    16'hCB85: data_out = 8'hD0;
                    16'hCB86: data_out = 8'hD1;
                    16'hCB87: data_out = 8'hD2;
                    16'hCB88: data_out = 8'hD3;
                    16'hCB89: data_out = 8'hD4;
                    16'hCB8A: data_out = 8'hD5;
                    16'hCB8B: data_out = 8'hD6;
                    16'hCB8C: data_out = 8'hD7;
                    16'hCB8D: data_out = 8'hD8;
                    16'hCB8E: data_out = 8'hD9;
                    16'hCB8F: data_out = 8'hDA;
                    16'hCB90: data_out = 8'hDB;
                    16'hCB91: data_out = 8'hDC;
                    16'hCB92: data_out = 8'hDD;
                    16'hCB93: data_out = 8'hDE;
                    16'hCB94: data_out = 8'hDF;
                    16'hCB95: data_out = 8'hE0;
                    16'hCB96: data_out = 8'hE1;
                    16'hCB97: data_out = 8'hE2;
                    16'hCB98: data_out = 8'hE3;
                    16'hCB99: data_out = 8'hE4;
                    16'hCB9A: data_out = 8'hE5;
                    16'hCB9B: data_out = 8'hE6;
                    16'hCB9C: data_out = 8'hE7;
                    16'hCB9D: data_out = 8'hE8;
                    16'hCB9E: data_out = 8'hE9;
                    16'hCB9F: data_out = 8'hEA;
                    16'hCBA0: data_out = 8'hEB;
                    16'hCBA1: data_out = 8'hEC;
                    16'hCBA2: data_out = 8'hED;
                    16'hCBA3: data_out = 8'hEE;
                    16'hCBA4: data_out = 8'hEF;
                    16'hCBA5: data_out = 8'hF0;
                    16'hCBA6: data_out = 8'hF1;
                    16'hCBA7: data_out = 8'hF2;
                    16'hCBA8: data_out = 8'hF3;
                    16'hCBA9: data_out = 8'hF4;
                    16'hCBAA: data_out = 8'hF5;
                    16'hCBAB: data_out = 8'hF6;
                    16'hCBAC: data_out = 8'hF7;
                    16'hCBAD: data_out = 8'hF8;
                    16'hCBAE: data_out = 8'hF9;
                    16'hCBAF: data_out = 8'hFA;
                    16'hCBB0: data_out = 8'hFB;
                    16'hCBB1: data_out = 8'hFC;
                    16'hCBB2: data_out = 8'hFD;
                    16'hCBB3: data_out = 8'hFE;
                    16'hCBB4: data_out = 8'hFF;
                    16'hCBB5: data_out = 8'h80;
                    16'hCBB6: data_out = 8'h81;
                    16'hCBB7: data_out = 8'h82;
                    16'hCBB8: data_out = 8'h83;
                    16'hCBB9: data_out = 8'h84;
                    16'hCBBA: data_out = 8'h85;
                    16'hCBBB: data_out = 8'h86;
                    16'hCBBC: data_out = 8'h87;
                    16'hCBBD: data_out = 8'h88;
                    16'hCBBE: data_out = 8'h89;
                    16'hCBBF: data_out = 8'h8A;
                    16'hCBC0: data_out = 8'h8B;
                    16'hCBC1: data_out = 8'h8C;
                    16'hCBC2: data_out = 8'h8D;
                    16'hCBC3: data_out = 8'h8E;
                    16'hCBC4: data_out = 8'h8F;
                    16'hCBC5: data_out = 8'h90;
                    16'hCBC6: data_out = 8'h91;
                    16'hCBC7: data_out = 8'h92;
                    16'hCBC8: data_out = 8'h93;
                    16'hCBC9: data_out = 8'h94;
                    16'hCBCA: data_out = 8'h95;
                    16'hCBCB: data_out = 8'h96;
                    16'hCBCC: data_out = 8'h97;
                    16'hCBCD: data_out = 8'h98;
                    16'hCBCE: data_out = 8'h99;
                    16'hCBCF: data_out = 8'h9A;
                    16'hCBD0: data_out = 8'h9B;
                    16'hCBD1: data_out = 8'h9C;
                    16'hCBD2: data_out = 8'h9D;
                    16'hCBD3: data_out = 8'h9E;
                    16'hCBD4: data_out = 8'h9F;
                    16'hCBD5: data_out = 8'hA0;
                    16'hCBD6: data_out = 8'hA1;
                    16'hCBD7: data_out = 8'hA2;
                    16'hCBD8: data_out = 8'hA3;
                    16'hCBD9: data_out = 8'hA4;
                    16'hCBDA: data_out = 8'hA5;
                    16'hCBDB: data_out = 8'hA6;
                    16'hCBDC: data_out = 8'hA7;
                    16'hCBDD: data_out = 8'hA8;
                    16'hCBDE: data_out = 8'hA9;
                    16'hCBDF: data_out = 8'hAA;
                    16'hCBE0: data_out = 8'hAB;
                    16'hCBE1: data_out = 8'hAC;
                    16'hCBE2: data_out = 8'hAD;
                    16'hCBE3: data_out = 8'hAE;
                    16'hCBE4: data_out = 8'hAF;
                    16'hCBE5: data_out = 8'hB0;
                    16'hCBE6: data_out = 8'hB1;
                    16'hCBE7: data_out = 8'hB2;
                    16'hCBE8: data_out = 8'hB3;
                    16'hCBE9: data_out = 8'hB4;
                    16'hCBEA: data_out = 8'hB5;
                    16'hCBEB: data_out = 8'hB6;
                    16'hCBEC: data_out = 8'hB7;
                    16'hCBED: data_out = 8'hB8;
                    16'hCBEE: data_out = 8'hB9;
                    16'hCBEF: data_out = 8'hBA;
                    16'hCBF0: data_out = 8'hBB;
                    16'hCBF1: data_out = 8'hBC;
                    16'hCBF2: data_out = 8'hBD;
                    16'hCBF3: data_out = 8'hBE;
                    16'hCBF4: data_out = 8'hBF;
                    16'hCBF5: data_out = 8'hC0;
                    16'hCBF6: data_out = 8'hC1;
                    16'hCBF7: data_out = 8'hC2;
                    16'hCBF8: data_out = 8'hC3;
                    16'hCBF9: data_out = 8'hC4;
                    16'hCBFA: data_out = 8'hC5;
                    16'hCBFB: data_out = 8'hC6;
                    16'hCBFC: data_out = 8'hC7;
                    16'hCBFD: data_out = 8'hC8;
                    16'hCBFE: data_out = 8'hC9;
                    16'hCBFF: data_out = 8'hCA;
                    16'hCC00: data_out = 8'hCC;
                    16'hCC01: data_out = 8'hCB;
                    16'hCC02: data_out = 8'hCA;
                    16'hCC03: data_out = 8'hC9;
                    16'hCC04: data_out = 8'hC8;
                    16'hCC05: data_out = 8'hC7;
                    16'hCC06: data_out = 8'hC6;
                    16'hCC07: data_out = 8'hC5;
                    16'hCC08: data_out = 8'hC4;
                    16'hCC09: data_out = 8'hC3;
                    16'hCC0A: data_out = 8'hC2;
                    16'hCC0B: data_out = 8'hC1;
                    16'hCC0C: data_out = 8'hC0;
                    16'hCC0D: data_out = 8'hBF;
                    16'hCC0E: data_out = 8'hBE;
                    16'hCC0F: data_out = 8'hBD;
                    16'hCC10: data_out = 8'hBC;
                    16'hCC11: data_out = 8'hBB;
                    16'hCC12: data_out = 8'hBA;
                    16'hCC13: data_out = 8'hB9;
                    16'hCC14: data_out = 8'hB8;
                    16'hCC15: data_out = 8'hB7;
                    16'hCC16: data_out = 8'hB6;
                    16'hCC17: data_out = 8'hB5;
                    16'hCC18: data_out = 8'hB4;
                    16'hCC19: data_out = 8'hB3;
                    16'hCC1A: data_out = 8'hB2;
                    16'hCC1B: data_out = 8'hB1;
                    16'hCC1C: data_out = 8'hB0;
                    16'hCC1D: data_out = 8'hAF;
                    16'hCC1E: data_out = 8'hAE;
                    16'hCC1F: data_out = 8'hAD;
                    16'hCC20: data_out = 8'hAC;
                    16'hCC21: data_out = 8'hAB;
                    16'hCC22: data_out = 8'hAA;
                    16'hCC23: data_out = 8'hA9;
                    16'hCC24: data_out = 8'hA8;
                    16'hCC25: data_out = 8'hA7;
                    16'hCC26: data_out = 8'hA6;
                    16'hCC27: data_out = 8'hA5;
                    16'hCC28: data_out = 8'hA4;
                    16'hCC29: data_out = 8'hA3;
                    16'hCC2A: data_out = 8'hA2;
                    16'hCC2B: data_out = 8'hA1;
                    16'hCC2C: data_out = 8'hA0;
                    16'hCC2D: data_out = 8'h9F;
                    16'hCC2E: data_out = 8'h9E;
                    16'hCC2F: data_out = 8'h9D;
                    16'hCC30: data_out = 8'h9C;
                    16'hCC31: data_out = 8'h9B;
                    16'hCC32: data_out = 8'h9A;
                    16'hCC33: data_out = 8'h99;
                    16'hCC34: data_out = 8'h98;
                    16'hCC35: data_out = 8'h97;
                    16'hCC36: data_out = 8'h96;
                    16'hCC37: data_out = 8'h95;
                    16'hCC38: data_out = 8'h94;
                    16'hCC39: data_out = 8'h93;
                    16'hCC3A: data_out = 8'h92;
                    16'hCC3B: data_out = 8'h91;
                    16'hCC3C: data_out = 8'h90;
                    16'hCC3D: data_out = 8'h8F;
                    16'hCC3E: data_out = 8'h8E;
                    16'hCC3F: data_out = 8'h8D;
                    16'hCC40: data_out = 8'h8C;
                    16'hCC41: data_out = 8'h8B;
                    16'hCC42: data_out = 8'h8A;
                    16'hCC43: data_out = 8'h89;
                    16'hCC44: data_out = 8'h88;
                    16'hCC45: data_out = 8'h87;
                    16'hCC46: data_out = 8'h86;
                    16'hCC47: data_out = 8'h85;
                    16'hCC48: data_out = 8'h84;
                    16'hCC49: data_out = 8'h83;
                    16'hCC4A: data_out = 8'h82;
                    16'hCC4B: data_out = 8'h81;
                    16'hCC4C: data_out = 8'h0;
                    16'hCC4D: data_out = 8'h1;
                    16'hCC4E: data_out = 8'h2;
                    16'hCC4F: data_out = 8'h3;
                    16'hCC50: data_out = 8'h4;
                    16'hCC51: data_out = 8'h5;
                    16'hCC52: data_out = 8'h6;
                    16'hCC53: data_out = 8'h7;
                    16'hCC54: data_out = 8'h8;
                    16'hCC55: data_out = 8'h9;
                    16'hCC56: data_out = 8'hA;
                    16'hCC57: data_out = 8'hB;
                    16'hCC58: data_out = 8'hC;
                    16'hCC59: data_out = 8'hD;
                    16'hCC5A: data_out = 8'hE;
                    16'hCC5B: data_out = 8'hF;
                    16'hCC5C: data_out = 8'h10;
                    16'hCC5D: data_out = 8'h11;
                    16'hCC5E: data_out = 8'h12;
                    16'hCC5F: data_out = 8'h13;
                    16'hCC60: data_out = 8'h14;
                    16'hCC61: data_out = 8'h15;
                    16'hCC62: data_out = 8'h16;
                    16'hCC63: data_out = 8'h17;
                    16'hCC64: data_out = 8'h18;
                    16'hCC65: data_out = 8'h19;
                    16'hCC66: data_out = 8'h1A;
                    16'hCC67: data_out = 8'h1B;
                    16'hCC68: data_out = 8'h1C;
                    16'hCC69: data_out = 8'h1D;
                    16'hCC6A: data_out = 8'h1E;
                    16'hCC6B: data_out = 8'h1F;
                    16'hCC6C: data_out = 8'h20;
                    16'hCC6D: data_out = 8'h21;
                    16'hCC6E: data_out = 8'h22;
                    16'hCC6F: data_out = 8'h23;
                    16'hCC70: data_out = 8'h24;
                    16'hCC71: data_out = 8'h25;
                    16'hCC72: data_out = 8'h26;
                    16'hCC73: data_out = 8'h27;
                    16'hCC74: data_out = 8'h28;
                    16'hCC75: data_out = 8'h29;
                    16'hCC76: data_out = 8'h2A;
                    16'hCC77: data_out = 8'h2B;
                    16'hCC78: data_out = 8'h2C;
                    16'hCC79: data_out = 8'h2D;
                    16'hCC7A: data_out = 8'h2E;
                    16'hCC7B: data_out = 8'h2F;
                    16'hCC7C: data_out = 8'h30;
                    16'hCC7D: data_out = 8'h31;
                    16'hCC7E: data_out = 8'h32;
                    16'hCC7F: data_out = 8'h33;
                    16'hCC80: data_out = 8'hCC;
                    16'hCC81: data_out = 8'hCD;
                    16'hCC82: data_out = 8'hCE;
                    16'hCC83: data_out = 8'hCF;
                    16'hCC84: data_out = 8'hD0;
                    16'hCC85: data_out = 8'hD1;
                    16'hCC86: data_out = 8'hD2;
                    16'hCC87: data_out = 8'hD3;
                    16'hCC88: data_out = 8'hD4;
                    16'hCC89: data_out = 8'hD5;
                    16'hCC8A: data_out = 8'hD6;
                    16'hCC8B: data_out = 8'hD7;
                    16'hCC8C: data_out = 8'hD8;
                    16'hCC8D: data_out = 8'hD9;
                    16'hCC8E: data_out = 8'hDA;
                    16'hCC8F: data_out = 8'hDB;
                    16'hCC90: data_out = 8'hDC;
                    16'hCC91: data_out = 8'hDD;
                    16'hCC92: data_out = 8'hDE;
                    16'hCC93: data_out = 8'hDF;
                    16'hCC94: data_out = 8'hE0;
                    16'hCC95: data_out = 8'hE1;
                    16'hCC96: data_out = 8'hE2;
                    16'hCC97: data_out = 8'hE3;
                    16'hCC98: data_out = 8'hE4;
                    16'hCC99: data_out = 8'hE5;
                    16'hCC9A: data_out = 8'hE6;
                    16'hCC9B: data_out = 8'hE7;
                    16'hCC9C: data_out = 8'hE8;
                    16'hCC9D: data_out = 8'hE9;
                    16'hCC9E: data_out = 8'hEA;
                    16'hCC9F: data_out = 8'hEB;
                    16'hCCA0: data_out = 8'hEC;
                    16'hCCA1: data_out = 8'hED;
                    16'hCCA2: data_out = 8'hEE;
                    16'hCCA3: data_out = 8'hEF;
                    16'hCCA4: data_out = 8'hF0;
                    16'hCCA5: data_out = 8'hF1;
                    16'hCCA6: data_out = 8'hF2;
                    16'hCCA7: data_out = 8'hF3;
                    16'hCCA8: data_out = 8'hF4;
                    16'hCCA9: data_out = 8'hF5;
                    16'hCCAA: data_out = 8'hF6;
                    16'hCCAB: data_out = 8'hF7;
                    16'hCCAC: data_out = 8'hF8;
                    16'hCCAD: data_out = 8'hF9;
                    16'hCCAE: data_out = 8'hFA;
                    16'hCCAF: data_out = 8'hFB;
                    16'hCCB0: data_out = 8'hFC;
                    16'hCCB1: data_out = 8'hFD;
                    16'hCCB2: data_out = 8'hFE;
                    16'hCCB3: data_out = 8'hFF;
                    16'hCCB4: data_out = 8'h80;
                    16'hCCB5: data_out = 8'h81;
                    16'hCCB6: data_out = 8'h82;
                    16'hCCB7: data_out = 8'h83;
                    16'hCCB8: data_out = 8'h84;
                    16'hCCB9: data_out = 8'h85;
                    16'hCCBA: data_out = 8'h86;
                    16'hCCBB: data_out = 8'h87;
                    16'hCCBC: data_out = 8'h88;
                    16'hCCBD: data_out = 8'h89;
                    16'hCCBE: data_out = 8'h8A;
                    16'hCCBF: data_out = 8'h8B;
                    16'hCCC0: data_out = 8'h8C;
                    16'hCCC1: data_out = 8'h8D;
                    16'hCCC2: data_out = 8'h8E;
                    16'hCCC3: data_out = 8'h8F;
                    16'hCCC4: data_out = 8'h90;
                    16'hCCC5: data_out = 8'h91;
                    16'hCCC6: data_out = 8'h92;
                    16'hCCC7: data_out = 8'h93;
                    16'hCCC8: data_out = 8'h94;
                    16'hCCC9: data_out = 8'h95;
                    16'hCCCA: data_out = 8'h96;
                    16'hCCCB: data_out = 8'h97;
                    16'hCCCC: data_out = 8'h98;
                    16'hCCCD: data_out = 8'h99;
                    16'hCCCE: data_out = 8'h9A;
                    16'hCCCF: data_out = 8'h9B;
                    16'hCCD0: data_out = 8'h9C;
                    16'hCCD1: data_out = 8'h9D;
                    16'hCCD2: data_out = 8'h9E;
                    16'hCCD3: data_out = 8'h9F;
                    16'hCCD4: data_out = 8'hA0;
                    16'hCCD5: data_out = 8'hA1;
                    16'hCCD6: data_out = 8'hA2;
                    16'hCCD7: data_out = 8'hA3;
                    16'hCCD8: data_out = 8'hA4;
                    16'hCCD9: data_out = 8'hA5;
                    16'hCCDA: data_out = 8'hA6;
                    16'hCCDB: data_out = 8'hA7;
                    16'hCCDC: data_out = 8'hA8;
                    16'hCCDD: data_out = 8'hA9;
                    16'hCCDE: data_out = 8'hAA;
                    16'hCCDF: data_out = 8'hAB;
                    16'hCCE0: data_out = 8'hAC;
                    16'hCCE1: data_out = 8'hAD;
                    16'hCCE2: data_out = 8'hAE;
                    16'hCCE3: data_out = 8'hAF;
                    16'hCCE4: data_out = 8'hB0;
                    16'hCCE5: data_out = 8'hB1;
                    16'hCCE6: data_out = 8'hB2;
                    16'hCCE7: data_out = 8'hB3;
                    16'hCCE8: data_out = 8'hB4;
                    16'hCCE9: data_out = 8'hB5;
                    16'hCCEA: data_out = 8'hB6;
                    16'hCCEB: data_out = 8'hB7;
                    16'hCCEC: data_out = 8'hB8;
                    16'hCCED: data_out = 8'hB9;
                    16'hCCEE: data_out = 8'hBA;
                    16'hCCEF: data_out = 8'hBB;
                    16'hCCF0: data_out = 8'hBC;
                    16'hCCF1: data_out = 8'hBD;
                    16'hCCF2: data_out = 8'hBE;
                    16'hCCF3: data_out = 8'hBF;
                    16'hCCF4: data_out = 8'hC0;
                    16'hCCF5: data_out = 8'hC1;
                    16'hCCF6: data_out = 8'hC2;
                    16'hCCF7: data_out = 8'hC3;
                    16'hCCF8: data_out = 8'hC4;
                    16'hCCF9: data_out = 8'hC5;
                    16'hCCFA: data_out = 8'hC6;
                    16'hCCFB: data_out = 8'hC7;
                    16'hCCFC: data_out = 8'hC8;
                    16'hCCFD: data_out = 8'hC9;
                    16'hCCFE: data_out = 8'hCA;
                    16'hCCFF: data_out = 8'hCB;
                    16'hCD00: data_out = 8'hCD;
                    16'hCD01: data_out = 8'hCC;
                    16'hCD02: data_out = 8'hCB;
                    16'hCD03: data_out = 8'hCA;
                    16'hCD04: data_out = 8'hC9;
                    16'hCD05: data_out = 8'hC8;
                    16'hCD06: data_out = 8'hC7;
                    16'hCD07: data_out = 8'hC6;
                    16'hCD08: data_out = 8'hC5;
                    16'hCD09: data_out = 8'hC4;
                    16'hCD0A: data_out = 8'hC3;
                    16'hCD0B: data_out = 8'hC2;
                    16'hCD0C: data_out = 8'hC1;
                    16'hCD0D: data_out = 8'hC0;
                    16'hCD0E: data_out = 8'hBF;
                    16'hCD0F: data_out = 8'hBE;
                    16'hCD10: data_out = 8'hBD;
                    16'hCD11: data_out = 8'hBC;
                    16'hCD12: data_out = 8'hBB;
                    16'hCD13: data_out = 8'hBA;
                    16'hCD14: data_out = 8'hB9;
                    16'hCD15: data_out = 8'hB8;
                    16'hCD16: data_out = 8'hB7;
                    16'hCD17: data_out = 8'hB6;
                    16'hCD18: data_out = 8'hB5;
                    16'hCD19: data_out = 8'hB4;
                    16'hCD1A: data_out = 8'hB3;
                    16'hCD1B: data_out = 8'hB2;
                    16'hCD1C: data_out = 8'hB1;
                    16'hCD1D: data_out = 8'hB0;
                    16'hCD1E: data_out = 8'hAF;
                    16'hCD1F: data_out = 8'hAE;
                    16'hCD20: data_out = 8'hAD;
                    16'hCD21: data_out = 8'hAC;
                    16'hCD22: data_out = 8'hAB;
                    16'hCD23: data_out = 8'hAA;
                    16'hCD24: data_out = 8'hA9;
                    16'hCD25: data_out = 8'hA8;
                    16'hCD26: data_out = 8'hA7;
                    16'hCD27: data_out = 8'hA6;
                    16'hCD28: data_out = 8'hA5;
                    16'hCD29: data_out = 8'hA4;
                    16'hCD2A: data_out = 8'hA3;
                    16'hCD2B: data_out = 8'hA2;
                    16'hCD2C: data_out = 8'hA1;
                    16'hCD2D: data_out = 8'hA0;
                    16'hCD2E: data_out = 8'h9F;
                    16'hCD2F: data_out = 8'h9E;
                    16'hCD30: data_out = 8'h9D;
                    16'hCD31: data_out = 8'h9C;
                    16'hCD32: data_out = 8'h9B;
                    16'hCD33: data_out = 8'h9A;
                    16'hCD34: data_out = 8'h99;
                    16'hCD35: data_out = 8'h98;
                    16'hCD36: data_out = 8'h97;
                    16'hCD37: data_out = 8'h96;
                    16'hCD38: data_out = 8'h95;
                    16'hCD39: data_out = 8'h94;
                    16'hCD3A: data_out = 8'h93;
                    16'hCD3B: data_out = 8'h92;
                    16'hCD3C: data_out = 8'h91;
                    16'hCD3D: data_out = 8'h90;
                    16'hCD3E: data_out = 8'h8F;
                    16'hCD3F: data_out = 8'h8E;
                    16'hCD40: data_out = 8'h8D;
                    16'hCD41: data_out = 8'h8C;
                    16'hCD42: data_out = 8'h8B;
                    16'hCD43: data_out = 8'h8A;
                    16'hCD44: data_out = 8'h89;
                    16'hCD45: data_out = 8'h88;
                    16'hCD46: data_out = 8'h87;
                    16'hCD47: data_out = 8'h86;
                    16'hCD48: data_out = 8'h85;
                    16'hCD49: data_out = 8'h84;
                    16'hCD4A: data_out = 8'h83;
                    16'hCD4B: data_out = 8'h82;
                    16'hCD4C: data_out = 8'h81;
                    16'hCD4D: data_out = 8'h0;
                    16'hCD4E: data_out = 8'h1;
                    16'hCD4F: data_out = 8'h2;
                    16'hCD50: data_out = 8'h3;
                    16'hCD51: data_out = 8'h4;
                    16'hCD52: data_out = 8'h5;
                    16'hCD53: data_out = 8'h6;
                    16'hCD54: data_out = 8'h7;
                    16'hCD55: data_out = 8'h8;
                    16'hCD56: data_out = 8'h9;
                    16'hCD57: data_out = 8'hA;
                    16'hCD58: data_out = 8'hB;
                    16'hCD59: data_out = 8'hC;
                    16'hCD5A: data_out = 8'hD;
                    16'hCD5B: data_out = 8'hE;
                    16'hCD5C: data_out = 8'hF;
                    16'hCD5D: data_out = 8'h10;
                    16'hCD5E: data_out = 8'h11;
                    16'hCD5F: data_out = 8'h12;
                    16'hCD60: data_out = 8'h13;
                    16'hCD61: data_out = 8'h14;
                    16'hCD62: data_out = 8'h15;
                    16'hCD63: data_out = 8'h16;
                    16'hCD64: data_out = 8'h17;
                    16'hCD65: data_out = 8'h18;
                    16'hCD66: data_out = 8'h19;
                    16'hCD67: data_out = 8'h1A;
                    16'hCD68: data_out = 8'h1B;
                    16'hCD69: data_out = 8'h1C;
                    16'hCD6A: data_out = 8'h1D;
                    16'hCD6B: data_out = 8'h1E;
                    16'hCD6C: data_out = 8'h1F;
                    16'hCD6D: data_out = 8'h20;
                    16'hCD6E: data_out = 8'h21;
                    16'hCD6F: data_out = 8'h22;
                    16'hCD70: data_out = 8'h23;
                    16'hCD71: data_out = 8'h24;
                    16'hCD72: data_out = 8'h25;
                    16'hCD73: data_out = 8'h26;
                    16'hCD74: data_out = 8'h27;
                    16'hCD75: data_out = 8'h28;
                    16'hCD76: data_out = 8'h29;
                    16'hCD77: data_out = 8'h2A;
                    16'hCD78: data_out = 8'h2B;
                    16'hCD79: data_out = 8'h2C;
                    16'hCD7A: data_out = 8'h2D;
                    16'hCD7B: data_out = 8'h2E;
                    16'hCD7C: data_out = 8'h2F;
                    16'hCD7D: data_out = 8'h30;
                    16'hCD7E: data_out = 8'h31;
                    16'hCD7F: data_out = 8'h32;
                    16'hCD80: data_out = 8'hCD;
                    16'hCD81: data_out = 8'hCE;
                    16'hCD82: data_out = 8'hCF;
                    16'hCD83: data_out = 8'hD0;
                    16'hCD84: data_out = 8'hD1;
                    16'hCD85: data_out = 8'hD2;
                    16'hCD86: data_out = 8'hD3;
                    16'hCD87: data_out = 8'hD4;
                    16'hCD88: data_out = 8'hD5;
                    16'hCD89: data_out = 8'hD6;
                    16'hCD8A: data_out = 8'hD7;
                    16'hCD8B: data_out = 8'hD8;
                    16'hCD8C: data_out = 8'hD9;
                    16'hCD8D: data_out = 8'hDA;
                    16'hCD8E: data_out = 8'hDB;
                    16'hCD8F: data_out = 8'hDC;
                    16'hCD90: data_out = 8'hDD;
                    16'hCD91: data_out = 8'hDE;
                    16'hCD92: data_out = 8'hDF;
                    16'hCD93: data_out = 8'hE0;
                    16'hCD94: data_out = 8'hE1;
                    16'hCD95: data_out = 8'hE2;
                    16'hCD96: data_out = 8'hE3;
                    16'hCD97: data_out = 8'hE4;
                    16'hCD98: data_out = 8'hE5;
                    16'hCD99: data_out = 8'hE6;
                    16'hCD9A: data_out = 8'hE7;
                    16'hCD9B: data_out = 8'hE8;
                    16'hCD9C: data_out = 8'hE9;
                    16'hCD9D: data_out = 8'hEA;
                    16'hCD9E: data_out = 8'hEB;
                    16'hCD9F: data_out = 8'hEC;
                    16'hCDA0: data_out = 8'hED;
                    16'hCDA1: data_out = 8'hEE;
                    16'hCDA2: data_out = 8'hEF;
                    16'hCDA3: data_out = 8'hF0;
                    16'hCDA4: data_out = 8'hF1;
                    16'hCDA5: data_out = 8'hF2;
                    16'hCDA6: data_out = 8'hF3;
                    16'hCDA7: data_out = 8'hF4;
                    16'hCDA8: data_out = 8'hF5;
                    16'hCDA9: data_out = 8'hF6;
                    16'hCDAA: data_out = 8'hF7;
                    16'hCDAB: data_out = 8'hF8;
                    16'hCDAC: data_out = 8'hF9;
                    16'hCDAD: data_out = 8'hFA;
                    16'hCDAE: data_out = 8'hFB;
                    16'hCDAF: data_out = 8'hFC;
                    16'hCDB0: data_out = 8'hFD;
                    16'hCDB1: data_out = 8'hFE;
                    16'hCDB2: data_out = 8'hFF;
                    16'hCDB3: data_out = 8'h80;
                    16'hCDB4: data_out = 8'h81;
                    16'hCDB5: data_out = 8'h82;
                    16'hCDB6: data_out = 8'h83;
                    16'hCDB7: data_out = 8'h84;
                    16'hCDB8: data_out = 8'h85;
                    16'hCDB9: data_out = 8'h86;
                    16'hCDBA: data_out = 8'h87;
                    16'hCDBB: data_out = 8'h88;
                    16'hCDBC: data_out = 8'h89;
                    16'hCDBD: data_out = 8'h8A;
                    16'hCDBE: data_out = 8'h8B;
                    16'hCDBF: data_out = 8'h8C;
                    16'hCDC0: data_out = 8'h8D;
                    16'hCDC1: data_out = 8'h8E;
                    16'hCDC2: data_out = 8'h8F;
                    16'hCDC3: data_out = 8'h90;
                    16'hCDC4: data_out = 8'h91;
                    16'hCDC5: data_out = 8'h92;
                    16'hCDC6: data_out = 8'h93;
                    16'hCDC7: data_out = 8'h94;
                    16'hCDC8: data_out = 8'h95;
                    16'hCDC9: data_out = 8'h96;
                    16'hCDCA: data_out = 8'h97;
                    16'hCDCB: data_out = 8'h98;
                    16'hCDCC: data_out = 8'h99;
                    16'hCDCD: data_out = 8'h9A;
                    16'hCDCE: data_out = 8'h9B;
                    16'hCDCF: data_out = 8'h9C;
                    16'hCDD0: data_out = 8'h9D;
                    16'hCDD1: data_out = 8'h9E;
                    16'hCDD2: data_out = 8'h9F;
                    16'hCDD3: data_out = 8'hA0;
                    16'hCDD4: data_out = 8'hA1;
                    16'hCDD5: data_out = 8'hA2;
                    16'hCDD6: data_out = 8'hA3;
                    16'hCDD7: data_out = 8'hA4;
                    16'hCDD8: data_out = 8'hA5;
                    16'hCDD9: data_out = 8'hA6;
                    16'hCDDA: data_out = 8'hA7;
                    16'hCDDB: data_out = 8'hA8;
                    16'hCDDC: data_out = 8'hA9;
                    16'hCDDD: data_out = 8'hAA;
                    16'hCDDE: data_out = 8'hAB;
                    16'hCDDF: data_out = 8'hAC;
                    16'hCDE0: data_out = 8'hAD;
                    16'hCDE1: data_out = 8'hAE;
                    16'hCDE2: data_out = 8'hAF;
                    16'hCDE3: data_out = 8'hB0;
                    16'hCDE4: data_out = 8'hB1;
                    16'hCDE5: data_out = 8'hB2;
                    16'hCDE6: data_out = 8'hB3;
                    16'hCDE7: data_out = 8'hB4;
                    16'hCDE8: data_out = 8'hB5;
                    16'hCDE9: data_out = 8'hB6;
                    16'hCDEA: data_out = 8'hB7;
                    16'hCDEB: data_out = 8'hB8;
                    16'hCDEC: data_out = 8'hB9;
                    16'hCDED: data_out = 8'hBA;
                    16'hCDEE: data_out = 8'hBB;
                    16'hCDEF: data_out = 8'hBC;
                    16'hCDF0: data_out = 8'hBD;
                    16'hCDF1: data_out = 8'hBE;
                    16'hCDF2: data_out = 8'hBF;
                    16'hCDF3: data_out = 8'hC0;
                    16'hCDF4: data_out = 8'hC1;
                    16'hCDF5: data_out = 8'hC2;
                    16'hCDF6: data_out = 8'hC3;
                    16'hCDF7: data_out = 8'hC4;
                    16'hCDF8: data_out = 8'hC5;
                    16'hCDF9: data_out = 8'hC6;
                    16'hCDFA: data_out = 8'hC7;
                    16'hCDFB: data_out = 8'hC8;
                    16'hCDFC: data_out = 8'hC9;
                    16'hCDFD: data_out = 8'hCA;
                    16'hCDFE: data_out = 8'hCB;
                    16'hCDFF: data_out = 8'hCC;
                    16'hCE00: data_out = 8'hCE;
                    16'hCE01: data_out = 8'hCD;
                    16'hCE02: data_out = 8'hCC;
                    16'hCE03: data_out = 8'hCB;
                    16'hCE04: data_out = 8'hCA;
                    16'hCE05: data_out = 8'hC9;
                    16'hCE06: data_out = 8'hC8;
                    16'hCE07: data_out = 8'hC7;
                    16'hCE08: data_out = 8'hC6;
                    16'hCE09: data_out = 8'hC5;
                    16'hCE0A: data_out = 8'hC4;
                    16'hCE0B: data_out = 8'hC3;
                    16'hCE0C: data_out = 8'hC2;
                    16'hCE0D: data_out = 8'hC1;
                    16'hCE0E: data_out = 8'hC0;
                    16'hCE0F: data_out = 8'hBF;
                    16'hCE10: data_out = 8'hBE;
                    16'hCE11: data_out = 8'hBD;
                    16'hCE12: data_out = 8'hBC;
                    16'hCE13: data_out = 8'hBB;
                    16'hCE14: data_out = 8'hBA;
                    16'hCE15: data_out = 8'hB9;
                    16'hCE16: data_out = 8'hB8;
                    16'hCE17: data_out = 8'hB7;
                    16'hCE18: data_out = 8'hB6;
                    16'hCE19: data_out = 8'hB5;
                    16'hCE1A: data_out = 8'hB4;
                    16'hCE1B: data_out = 8'hB3;
                    16'hCE1C: data_out = 8'hB2;
                    16'hCE1D: data_out = 8'hB1;
                    16'hCE1E: data_out = 8'hB0;
                    16'hCE1F: data_out = 8'hAF;
                    16'hCE20: data_out = 8'hAE;
                    16'hCE21: data_out = 8'hAD;
                    16'hCE22: data_out = 8'hAC;
                    16'hCE23: data_out = 8'hAB;
                    16'hCE24: data_out = 8'hAA;
                    16'hCE25: data_out = 8'hA9;
                    16'hCE26: data_out = 8'hA8;
                    16'hCE27: data_out = 8'hA7;
                    16'hCE28: data_out = 8'hA6;
                    16'hCE29: data_out = 8'hA5;
                    16'hCE2A: data_out = 8'hA4;
                    16'hCE2B: data_out = 8'hA3;
                    16'hCE2C: data_out = 8'hA2;
                    16'hCE2D: data_out = 8'hA1;
                    16'hCE2E: data_out = 8'hA0;
                    16'hCE2F: data_out = 8'h9F;
                    16'hCE30: data_out = 8'h9E;
                    16'hCE31: data_out = 8'h9D;
                    16'hCE32: data_out = 8'h9C;
                    16'hCE33: data_out = 8'h9B;
                    16'hCE34: data_out = 8'h9A;
                    16'hCE35: data_out = 8'h99;
                    16'hCE36: data_out = 8'h98;
                    16'hCE37: data_out = 8'h97;
                    16'hCE38: data_out = 8'h96;
                    16'hCE39: data_out = 8'h95;
                    16'hCE3A: data_out = 8'h94;
                    16'hCE3B: data_out = 8'h93;
                    16'hCE3C: data_out = 8'h92;
                    16'hCE3D: data_out = 8'h91;
                    16'hCE3E: data_out = 8'h90;
                    16'hCE3F: data_out = 8'h8F;
                    16'hCE40: data_out = 8'h8E;
                    16'hCE41: data_out = 8'h8D;
                    16'hCE42: data_out = 8'h8C;
                    16'hCE43: data_out = 8'h8B;
                    16'hCE44: data_out = 8'h8A;
                    16'hCE45: data_out = 8'h89;
                    16'hCE46: data_out = 8'h88;
                    16'hCE47: data_out = 8'h87;
                    16'hCE48: data_out = 8'h86;
                    16'hCE49: data_out = 8'h85;
                    16'hCE4A: data_out = 8'h84;
                    16'hCE4B: data_out = 8'h83;
                    16'hCE4C: data_out = 8'h82;
                    16'hCE4D: data_out = 8'h81;
                    16'hCE4E: data_out = 8'h0;
                    16'hCE4F: data_out = 8'h1;
                    16'hCE50: data_out = 8'h2;
                    16'hCE51: data_out = 8'h3;
                    16'hCE52: data_out = 8'h4;
                    16'hCE53: data_out = 8'h5;
                    16'hCE54: data_out = 8'h6;
                    16'hCE55: data_out = 8'h7;
                    16'hCE56: data_out = 8'h8;
                    16'hCE57: data_out = 8'h9;
                    16'hCE58: data_out = 8'hA;
                    16'hCE59: data_out = 8'hB;
                    16'hCE5A: data_out = 8'hC;
                    16'hCE5B: data_out = 8'hD;
                    16'hCE5C: data_out = 8'hE;
                    16'hCE5D: data_out = 8'hF;
                    16'hCE5E: data_out = 8'h10;
                    16'hCE5F: data_out = 8'h11;
                    16'hCE60: data_out = 8'h12;
                    16'hCE61: data_out = 8'h13;
                    16'hCE62: data_out = 8'h14;
                    16'hCE63: data_out = 8'h15;
                    16'hCE64: data_out = 8'h16;
                    16'hCE65: data_out = 8'h17;
                    16'hCE66: data_out = 8'h18;
                    16'hCE67: data_out = 8'h19;
                    16'hCE68: data_out = 8'h1A;
                    16'hCE69: data_out = 8'h1B;
                    16'hCE6A: data_out = 8'h1C;
                    16'hCE6B: data_out = 8'h1D;
                    16'hCE6C: data_out = 8'h1E;
                    16'hCE6D: data_out = 8'h1F;
                    16'hCE6E: data_out = 8'h20;
                    16'hCE6F: data_out = 8'h21;
                    16'hCE70: data_out = 8'h22;
                    16'hCE71: data_out = 8'h23;
                    16'hCE72: data_out = 8'h24;
                    16'hCE73: data_out = 8'h25;
                    16'hCE74: data_out = 8'h26;
                    16'hCE75: data_out = 8'h27;
                    16'hCE76: data_out = 8'h28;
                    16'hCE77: data_out = 8'h29;
                    16'hCE78: data_out = 8'h2A;
                    16'hCE79: data_out = 8'h2B;
                    16'hCE7A: data_out = 8'h2C;
                    16'hCE7B: data_out = 8'h2D;
                    16'hCE7C: data_out = 8'h2E;
                    16'hCE7D: data_out = 8'h2F;
                    16'hCE7E: data_out = 8'h30;
                    16'hCE7F: data_out = 8'h31;
                    16'hCE80: data_out = 8'hCE;
                    16'hCE81: data_out = 8'hCF;
                    16'hCE82: data_out = 8'hD0;
                    16'hCE83: data_out = 8'hD1;
                    16'hCE84: data_out = 8'hD2;
                    16'hCE85: data_out = 8'hD3;
                    16'hCE86: data_out = 8'hD4;
                    16'hCE87: data_out = 8'hD5;
                    16'hCE88: data_out = 8'hD6;
                    16'hCE89: data_out = 8'hD7;
                    16'hCE8A: data_out = 8'hD8;
                    16'hCE8B: data_out = 8'hD9;
                    16'hCE8C: data_out = 8'hDA;
                    16'hCE8D: data_out = 8'hDB;
                    16'hCE8E: data_out = 8'hDC;
                    16'hCE8F: data_out = 8'hDD;
                    16'hCE90: data_out = 8'hDE;
                    16'hCE91: data_out = 8'hDF;
                    16'hCE92: data_out = 8'hE0;
                    16'hCE93: data_out = 8'hE1;
                    16'hCE94: data_out = 8'hE2;
                    16'hCE95: data_out = 8'hE3;
                    16'hCE96: data_out = 8'hE4;
                    16'hCE97: data_out = 8'hE5;
                    16'hCE98: data_out = 8'hE6;
                    16'hCE99: data_out = 8'hE7;
                    16'hCE9A: data_out = 8'hE8;
                    16'hCE9B: data_out = 8'hE9;
                    16'hCE9C: data_out = 8'hEA;
                    16'hCE9D: data_out = 8'hEB;
                    16'hCE9E: data_out = 8'hEC;
                    16'hCE9F: data_out = 8'hED;
                    16'hCEA0: data_out = 8'hEE;
                    16'hCEA1: data_out = 8'hEF;
                    16'hCEA2: data_out = 8'hF0;
                    16'hCEA3: data_out = 8'hF1;
                    16'hCEA4: data_out = 8'hF2;
                    16'hCEA5: data_out = 8'hF3;
                    16'hCEA6: data_out = 8'hF4;
                    16'hCEA7: data_out = 8'hF5;
                    16'hCEA8: data_out = 8'hF6;
                    16'hCEA9: data_out = 8'hF7;
                    16'hCEAA: data_out = 8'hF8;
                    16'hCEAB: data_out = 8'hF9;
                    16'hCEAC: data_out = 8'hFA;
                    16'hCEAD: data_out = 8'hFB;
                    16'hCEAE: data_out = 8'hFC;
                    16'hCEAF: data_out = 8'hFD;
                    16'hCEB0: data_out = 8'hFE;
                    16'hCEB1: data_out = 8'hFF;
                    16'hCEB2: data_out = 8'h80;
                    16'hCEB3: data_out = 8'h81;
                    16'hCEB4: data_out = 8'h82;
                    16'hCEB5: data_out = 8'h83;
                    16'hCEB6: data_out = 8'h84;
                    16'hCEB7: data_out = 8'h85;
                    16'hCEB8: data_out = 8'h86;
                    16'hCEB9: data_out = 8'h87;
                    16'hCEBA: data_out = 8'h88;
                    16'hCEBB: data_out = 8'h89;
                    16'hCEBC: data_out = 8'h8A;
                    16'hCEBD: data_out = 8'h8B;
                    16'hCEBE: data_out = 8'h8C;
                    16'hCEBF: data_out = 8'h8D;
                    16'hCEC0: data_out = 8'h8E;
                    16'hCEC1: data_out = 8'h8F;
                    16'hCEC2: data_out = 8'h90;
                    16'hCEC3: data_out = 8'h91;
                    16'hCEC4: data_out = 8'h92;
                    16'hCEC5: data_out = 8'h93;
                    16'hCEC6: data_out = 8'h94;
                    16'hCEC7: data_out = 8'h95;
                    16'hCEC8: data_out = 8'h96;
                    16'hCEC9: data_out = 8'h97;
                    16'hCECA: data_out = 8'h98;
                    16'hCECB: data_out = 8'h99;
                    16'hCECC: data_out = 8'h9A;
                    16'hCECD: data_out = 8'h9B;
                    16'hCECE: data_out = 8'h9C;
                    16'hCECF: data_out = 8'h9D;
                    16'hCED0: data_out = 8'h9E;
                    16'hCED1: data_out = 8'h9F;
                    16'hCED2: data_out = 8'hA0;
                    16'hCED3: data_out = 8'hA1;
                    16'hCED4: data_out = 8'hA2;
                    16'hCED5: data_out = 8'hA3;
                    16'hCED6: data_out = 8'hA4;
                    16'hCED7: data_out = 8'hA5;
                    16'hCED8: data_out = 8'hA6;
                    16'hCED9: data_out = 8'hA7;
                    16'hCEDA: data_out = 8'hA8;
                    16'hCEDB: data_out = 8'hA9;
                    16'hCEDC: data_out = 8'hAA;
                    16'hCEDD: data_out = 8'hAB;
                    16'hCEDE: data_out = 8'hAC;
                    16'hCEDF: data_out = 8'hAD;
                    16'hCEE0: data_out = 8'hAE;
                    16'hCEE1: data_out = 8'hAF;
                    16'hCEE2: data_out = 8'hB0;
                    16'hCEE3: data_out = 8'hB1;
                    16'hCEE4: data_out = 8'hB2;
                    16'hCEE5: data_out = 8'hB3;
                    16'hCEE6: data_out = 8'hB4;
                    16'hCEE7: data_out = 8'hB5;
                    16'hCEE8: data_out = 8'hB6;
                    16'hCEE9: data_out = 8'hB7;
                    16'hCEEA: data_out = 8'hB8;
                    16'hCEEB: data_out = 8'hB9;
                    16'hCEEC: data_out = 8'hBA;
                    16'hCEED: data_out = 8'hBB;
                    16'hCEEE: data_out = 8'hBC;
                    16'hCEEF: data_out = 8'hBD;
                    16'hCEF0: data_out = 8'hBE;
                    16'hCEF1: data_out = 8'hBF;
                    16'hCEF2: data_out = 8'hC0;
                    16'hCEF3: data_out = 8'hC1;
                    16'hCEF4: data_out = 8'hC2;
                    16'hCEF5: data_out = 8'hC3;
                    16'hCEF6: data_out = 8'hC4;
                    16'hCEF7: data_out = 8'hC5;
                    16'hCEF8: data_out = 8'hC6;
                    16'hCEF9: data_out = 8'hC7;
                    16'hCEFA: data_out = 8'hC8;
                    16'hCEFB: data_out = 8'hC9;
                    16'hCEFC: data_out = 8'hCA;
                    16'hCEFD: data_out = 8'hCB;
                    16'hCEFE: data_out = 8'hCC;
                    16'hCEFF: data_out = 8'hCD;
                    16'hCF00: data_out = 8'hCF;
                    16'hCF01: data_out = 8'hCE;
                    16'hCF02: data_out = 8'hCD;
                    16'hCF03: data_out = 8'hCC;
                    16'hCF04: data_out = 8'hCB;
                    16'hCF05: data_out = 8'hCA;
                    16'hCF06: data_out = 8'hC9;
                    16'hCF07: data_out = 8'hC8;
                    16'hCF08: data_out = 8'hC7;
                    16'hCF09: data_out = 8'hC6;
                    16'hCF0A: data_out = 8'hC5;
                    16'hCF0B: data_out = 8'hC4;
                    16'hCF0C: data_out = 8'hC3;
                    16'hCF0D: data_out = 8'hC2;
                    16'hCF0E: data_out = 8'hC1;
                    16'hCF0F: data_out = 8'hC0;
                    16'hCF10: data_out = 8'hBF;
                    16'hCF11: data_out = 8'hBE;
                    16'hCF12: data_out = 8'hBD;
                    16'hCF13: data_out = 8'hBC;
                    16'hCF14: data_out = 8'hBB;
                    16'hCF15: data_out = 8'hBA;
                    16'hCF16: data_out = 8'hB9;
                    16'hCF17: data_out = 8'hB8;
                    16'hCF18: data_out = 8'hB7;
                    16'hCF19: data_out = 8'hB6;
                    16'hCF1A: data_out = 8'hB5;
                    16'hCF1B: data_out = 8'hB4;
                    16'hCF1C: data_out = 8'hB3;
                    16'hCF1D: data_out = 8'hB2;
                    16'hCF1E: data_out = 8'hB1;
                    16'hCF1F: data_out = 8'hB0;
                    16'hCF20: data_out = 8'hAF;
                    16'hCF21: data_out = 8'hAE;
                    16'hCF22: data_out = 8'hAD;
                    16'hCF23: data_out = 8'hAC;
                    16'hCF24: data_out = 8'hAB;
                    16'hCF25: data_out = 8'hAA;
                    16'hCF26: data_out = 8'hA9;
                    16'hCF27: data_out = 8'hA8;
                    16'hCF28: data_out = 8'hA7;
                    16'hCF29: data_out = 8'hA6;
                    16'hCF2A: data_out = 8'hA5;
                    16'hCF2B: data_out = 8'hA4;
                    16'hCF2C: data_out = 8'hA3;
                    16'hCF2D: data_out = 8'hA2;
                    16'hCF2E: data_out = 8'hA1;
                    16'hCF2F: data_out = 8'hA0;
                    16'hCF30: data_out = 8'h9F;
                    16'hCF31: data_out = 8'h9E;
                    16'hCF32: data_out = 8'h9D;
                    16'hCF33: data_out = 8'h9C;
                    16'hCF34: data_out = 8'h9B;
                    16'hCF35: data_out = 8'h9A;
                    16'hCF36: data_out = 8'h99;
                    16'hCF37: data_out = 8'h98;
                    16'hCF38: data_out = 8'h97;
                    16'hCF39: data_out = 8'h96;
                    16'hCF3A: data_out = 8'h95;
                    16'hCF3B: data_out = 8'h94;
                    16'hCF3C: data_out = 8'h93;
                    16'hCF3D: data_out = 8'h92;
                    16'hCF3E: data_out = 8'h91;
                    16'hCF3F: data_out = 8'h90;
                    16'hCF40: data_out = 8'h8F;
                    16'hCF41: data_out = 8'h8E;
                    16'hCF42: data_out = 8'h8D;
                    16'hCF43: data_out = 8'h8C;
                    16'hCF44: data_out = 8'h8B;
                    16'hCF45: data_out = 8'h8A;
                    16'hCF46: data_out = 8'h89;
                    16'hCF47: data_out = 8'h88;
                    16'hCF48: data_out = 8'h87;
                    16'hCF49: data_out = 8'h86;
                    16'hCF4A: data_out = 8'h85;
                    16'hCF4B: data_out = 8'h84;
                    16'hCF4C: data_out = 8'h83;
                    16'hCF4D: data_out = 8'h82;
                    16'hCF4E: data_out = 8'h81;
                    16'hCF4F: data_out = 8'h0;
                    16'hCF50: data_out = 8'h1;
                    16'hCF51: data_out = 8'h2;
                    16'hCF52: data_out = 8'h3;
                    16'hCF53: data_out = 8'h4;
                    16'hCF54: data_out = 8'h5;
                    16'hCF55: data_out = 8'h6;
                    16'hCF56: data_out = 8'h7;
                    16'hCF57: data_out = 8'h8;
                    16'hCF58: data_out = 8'h9;
                    16'hCF59: data_out = 8'hA;
                    16'hCF5A: data_out = 8'hB;
                    16'hCF5B: data_out = 8'hC;
                    16'hCF5C: data_out = 8'hD;
                    16'hCF5D: data_out = 8'hE;
                    16'hCF5E: data_out = 8'hF;
                    16'hCF5F: data_out = 8'h10;
                    16'hCF60: data_out = 8'h11;
                    16'hCF61: data_out = 8'h12;
                    16'hCF62: data_out = 8'h13;
                    16'hCF63: data_out = 8'h14;
                    16'hCF64: data_out = 8'h15;
                    16'hCF65: data_out = 8'h16;
                    16'hCF66: data_out = 8'h17;
                    16'hCF67: data_out = 8'h18;
                    16'hCF68: data_out = 8'h19;
                    16'hCF69: data_out = 8'h1A;
                    16'hCF6A: data_out = 8'h1B;
                    16'hCF6B: data_out = 8'h1C;
                    16'hCF6C: data_out = 8'h1D;
                    16'hCF6D: data_out = 8'h1E;
                    16'hCF6E: data_out = 8'h1F;
                    16'hCF6F: data_out = 8'h20;
                    16'hCF70: data_out = 8'h21;
                    16'hCF71: data_out = 8'h22;
                    16'hCF72: data_out = 8'h23;
                    16'hCF73: data_out = 8'h24;
                    16'hCF74: data_out = 8'h25;
                    16'hCF75: data_out = 8'h26;
                    16'hCF76: data_out = 8'h27;
                    16'hCF77: data_out = 8'h28;
                    16'hCF78: data_out = 8'h29;
                    16'hCF79: data_out = 8'h2A;
                    16'hCF7A: data_out = 8'h2B;
                    16'hCF7B: data_out = 8'h2C;
                    16'hCF7C: data_out = 8'h2D;
                    16'hCF7D: data_out = 8'h2E;
                    16'hCF7E: data_out = 8'h2F;
                    16'hCF7F: data_out = 8'h30;
                    16'hCF80: data_out = 8'hCF;
                    16'hCF81: data_out = 8'hD0;
                    16'hCF82: data_out = 8'hD1;
                    16'hCF83: data_out = 8'hD2;
                    16'hCF84: data_out = 8'hD3;
                    16'hCF85: data_out = 8'hD4;
                    16'hCF86: data_out = 8'hD5;
                    16'hCF87: data_out = 8'hD6;
                    16'hCF88: data_out = 8'hD7;
                    16'hCF89: data_out = 8'hD8;
                    16'hCF8A: data_out = 8'hD9;
                    16'hCF8B: data_out = 8'hDA;
                    16'hCF8C: data_out = 8'hDB;
                    16'hCF8D: data_out = 8'hDC;
                    16'hCF8E: data_out = 8'hDD;
                    16'hCF8F: data_out = 8'hDE;
                    16'hCF90: data_out = 8'hDF;
                    16'hCF91: data_out = 8'hE0;
                    16'hCF92: data_out = 8'hE1;
                    16'hCF93: data_out = 8'hE2;
                    16'hCF94: data_out = 8'hE3;
                    16'hCF95: data_out = 8'hE4;
                    16'hCF96: data_out = 8'hE5;
                    16'hCF97: data_out = 8'hE6;
                    16'hCF98: data_out = 8'hE7;
                    16'hCF99: data_out = 8'hE8;
                    16'hCF9A: data_out = 8'hE9;
                    16'hCF9B: data_out = 8'hEA;
                    16'hCF9C: data_out = 8'hEB;
                    16'hCF9D: data_out = 8'hEC;
                    16'hCF9E: data_out = 8'hED;
                    16'hCF9F: data_out = 8'hEE;
                    16'hCFA0: data_out = 8'hEF;
                    16'hCFA1: data_out = 8'hF0;
                    16'hCFA2: data_out = 8'hF1;
                    16'hCFA3: data_out = 8'hF2;
                    16'hCFA4: data_out = 8'hF3;
                    16'hCFA5: data_out = 8'hF4;
                    16'hCFA6: data_out = 8'hF5;
                    16'hCFA7: data_out = 8'hF6;
                    16'hCFA8: data_out = 8'hF7;
                    16'hCFA9: data_out = 8'hF8;
                    16'hCFAA: data_out = 8'hF9;
                    16'hCFAB: data_out = 8'hFA;
                    16'hCFAC: data_out = 8'hFB;
                    16'hCFAD: data_out = 8'hFC;
                    16'hCFAE: data_out = 8'hFD;
                    16'hCFAF: data_out = 8'hFE;
                    16'hCFB0: data_out = 8'hFF;
                    16'hCFB1: data_out = 8'h80;
                    16'hCFB2: data_out = 8'h81;
                    16'hCFB3: data_out = 8'h82;
                    16'hCFB4: data_out = 8'h83;
                    16'hCFB5: data_out = 8'h84;
                    16'hCFB6: data_out = 8'h85;
                    16'hCFB7: data_out = 8'h86;
                    16'hCFB8: data_out = 8'h87;
                    16'hCFB9: data_out = 8'h88;
                    16'hCFBA: data_out = 8'h89;
                    16'hCFBB: data_out = 8'h8A;
                    16'hCFBC: data_out = 8'h8B;
                    16'hCFBD: data_out = 8'h8C;
                    16'hCFBE: data_out = 8'h8D;
                    16'hCFBF: data_out = 8'h8E;
                    16'hCFC0: data_out = 8'h8F;
                    16'hCFC1: data_out = 8'h90;
                    16'hCFC2: data_out = 8'h91;
                    16'hCFC3: data_out = 8'h92;
                    16'hCFC4: data_out = 8'h93;
                    16'hCFC5: data_out = 8'h94;
                    16'hCFC6: data_out = 8'h95;
                    16'hCFC7: data_out = 8'h96;
                    16'hCFC8: data_out = 8'h97;
                    16'hCFC9: data_out = 8'h98;
                    16'hCFCA: data_out = 8'h99;
                    16'hCFCB: data_out = 8'h9A;
                    16'hCFCC: data_out = 8'h9B;
                    16'hCFCD: data_out = 8'h9C;
                    16'hCFCE: data_out = 8'h9D;
                    16'hCFCF: data_out = 8'h9E;
                    16'hCFD0: data_out = 8'h9F;
                    16'hCFD1: data_out = 8'hA0;
                    16'hCFD2: data_out = 8'hA1;
                    16'hCFD3: data_out = 8'hA2;
                    16'hCFD4: data_out = 8'hA3;
                    16'hCFD5: data_out = 8'hA4;
                    16'hCFD6: data_out = 8'hA5;
                    16'hCFD7: data_out = 8'hA6;
                    16'hCFD8: data_out = 8'hA7;
                    16'hCFD9: data_out = 8'hA8;
                    16'hCFDA: data_out = 8'hA9;
                    16'hCFDB: data_out = 8'hAA;
                    16'hCFDC: data_out = 8'hAB;
                    16'hCFDD: data_out = 8'hAC;
                    16'hCFDE: data_out = 8'hAD;
                    16'hCFDF: data_out = 8'hAE;
                    16'hCFE0: data_out = 8'hAF;
                    16'hCFE1: data_out = 8'hB0;
                    16'hCFE2: data_out = 8'hB1;
                    16'hCFE3: data_out = 8'hB2;
                    16'hCFE4: data_out = 8'hB3;
                    16'hCFE5: data_out = 8'hB4;
                    16'hCFE6: data_out = 8'hB5;
                    16'hCFE7: data_out = 8'hB6;
                    16'hCFE8: data_out = 8'hB7;
                    16'hCFE9: data_out = 8'hB8;
                    16'hCFEA: data_out = 8'hB9;
                    16'hCFEB: data_out = 8'hBA;
                    16'hCFEC: data_out = 8'hBB;
                    16'hCFED: data_out = 8'hBC;
                    16'hCFEE: data_out = 8'hBD;
                    16'hCFEF: data_out = 8'hBE;
                    16'hCFF0: data_out = 8'hBF;
                    16'hCFF1: data_out = 8'hC0;
                    16'hCFF2: data_out = 8'hC1;
                    16'hCFF3: data_out = 8'hC2;
                    16'hCFF4: data_out = 8'hC3;
                    16'hCFF5: data_out = 8'hC4;
                    16'hCFF6: data_out = 8'hC5;
                    16'hCFF7: data_out = 8'hC6;
                    16'hCFF8: data_out = 8'hC7;
                    16'hCFF9: data_out = 8'hC8;
                    16'hCFFA: data_out = 8'hC9;
                    16'hCFFB: data_out = 8'hCA;
                    16'hCFFC: data_out = 8'hCB;
                    16'hCFFD: data_out = 8'hCC;
                    16'hCFFE: data_out = 8'hCD;
                    16'hCFFF: data_out = 8'hCE;
                    16'hD000: data_out = 8'hD0;
                    16'hD001: data_out = 8'hCF;
                    16'hD002: data_out = 8'hCE;
                    16'hD003: data_out = 8'hCD;
                    16'hD004: data_out = 8'hCC;
                    16'hD005: data_out = 8'hCB;
                    16'hD006: data_out = 8'hCA;
                    16'hD007: data_out = 8'hC9;
                    16'hD008: data_out = 8'hC8;
                    16'hD009: data_out = 8'hC7;
                    16'hD00A: data_out = 8'hC6;
                    16'hD00B: data_out = 8'hC5;
                    16'hD00C: data_out = 8'hC4;
                    16'hD00D: data_out = 8'hC3;
                    16'hD00E: data_out = 8'hC2;
                    16'hD00F: data_out = 8'hC1;
                    16'hD010: data_out = 8'hC0;
                    16'hD011: data_out = 8'hBF;
                    16'hD012: data_out = 8'hBE;
                    16'hD013: data_out = 8'hBD;
                    16'hD014: data_out = 8'hBC;
                    16'hD015: data_out = 8'hBB;
                    16'hD016: data_out = 8'hBA;
                    16'hD017: data_out = 8'hB9;
                    16'hD018: data_out = 8'hB8;
                    16'hD019: data_out = 8'hB7;
                    16'hD01A: data_out = 8'hB6;
                    16'hD01B: data_out = 8'hB5;
                    16'hD01C: data_out = 8'hB4;
                    16'hD01D: data_out = 8'hB3;
                    16'hD01E: data_out = 8'hB2;
                    16'hD01F: data_out = 8'hB1;
                    16'hD020: data_out = 8'hB0;
                    16'hD021: data_out = 8'hAF;
                    16'hD022: data_out = 8'hAE;
                    16'hD023: data_out = 8'hAD;
                    16'hD024: data_out = 8'hAC;
                    16'hD025: data_out = 8'hAB;
                    16'hD026: data_out = 8'hAA;
                    16'hD027: data_out = 8'hA9;
                    16'hD028: data_out = 8'hA8;
                    16'hD029: data_out = 8'hA7;
                    16'hD02A: data_out = 8'hA6;
                    16'hD02B: data_out = 8'hA5;
                    16'hD02C: data_out = 8'hA4;
                    16'hD02D: data_out = 8'hA3;
                    16'hD02E: data_out = 8'hA2;
                    16'hD02F: data_out = 8'hA1;
                    16'hD030: data_out = 8'hA0;
                    16'hD031: data_out = 8'h9F;
                    16'hD032: data_out = 8'h9E;
                    16'hD033: data_out = 8'h9D;
                    16'hD034: data_out = 8'h9C;
                    16'hD035: data_out = 8'h9B;
                    16'hD036: data_out = 8'h9A;
                    16'hD037: data_out = 8'h99;
                    16'hD038: data_out = 8'h98;
                    16'hD039: data_out = 8'h97;
                    16'hD03A: data_out = 8'h96;
                    16'hD03B: data_out = 8'h95;
                    16'hD03C: data_out = 8'h94;
                    16'hD03D: data_out = 8'h93;
                    16'hD03E: data_out = 8'h92;
                    16'hD03F: data_out = 8'h91;
                    16'hD040: data_out = 8'h90;
                    16'hD041: data_out = 8'h8F;
                    16'hD042: data_out = 8'h8E;
                    16'hD043: data_out = 8'h8D;
                    16'hD044: data_out = 8'h8C;
                    16'hD045: data_out = 8'h8B;
                    16'hD046: data_out = 8'h8A;
                    16'hD047: data_out = 8'h89;
                    16'hD048: data_out = 8'h88;
                    16'hD049: data_out = 8'h87;
                    16'hD04A: data_out = 8'h86;
                    16'hD04B: data_out = 8'h85;
                    16'hD04C: data_out = 8'h84;
                    16'hD04D: data_out = 8'h83;
                    16'hD04E: data_out = 8'h82;
                    16'hD04F: data_out = 8'h81;
                    16'hD050: data_out = 8'h0;
                    16'hD051: data_out = 8'h1;
                    16'hD052: data_out = 8'h2;
                    16'hD053: data_out = 8'h3;
                    16'hD054: data_out = 8'h4;
                    16'hD055: data_out = 8'h5;
                    16'hD056: data_out = 8'h6;
                    16'hD057: data_out = 8'h7;
                    16'hD058: data_out = 8'h8;
                    16'hD059: data_out = 8'h9;
                    16'hD05A: data_out = 8'hA;
                    16'hD05B: data_out = 8'hB;
                    16'hD05C: data_out = 8'hC;
                    16'hD05D: data_out = 8'hD;
                    16'hD05E: data_out = 8'hE;
                    16'hD05F: data_out = 8'hF;
                    16'hD060: data_out = 8'h10;
                    16'hD061: data_out = 8'h11;
                    16'hD062: data_out = 8'h12;
                    16'hD063: data_out = 8'h13;
                    16'hD064: data_out = 8'h14;
                    16'hD065: data_out = 8'h15;
                    16'hD066: data_out = 8'h16;
                    16'hD067: data_out = 8'h17;
                    16'hD068: data_out = 8'h18;
                    16'hD069: data_out = 8'h19;
                    16'hD06A: data_out = 8'h1A;
                    16'hD06B: data_out = 8'h1B;
                    16'hD06C: data_out = 8'h1C;
                    16'hD06D: data_out = 8'h1D;
                    16'hD06E: data_out = 8'h1E;
                    16'hD06F: data_out = 8'h1F;
                    16'hD070: data_out = 8'h20;
                    16'hD071: data_out = 8'h21;
                    16'hD072: data_out = 8'h22;
                    16'hD073: data_out = 8'h23;
                    16'hD074: data_out = 8'h24;
                    16'hD075: data_out = 8'h25;
                    16'hD076: data_out = 8'h26;
                    16'hD077: data_out = 8'h27;
                    16'hD078: data_out = 8'h28;
                    16'hD079: data_out = 8'h29;
                    16'hD07A: data_out = 8'h2A;
                    16'hD07B: data_out = 8'h2B;
                    16'hD07C: data_out = 8'h2C;
                    16'hD07D: data_out = 8'h2D;
                    16'hD07E: data_out = 8'h2E;
                    16'hD07F: data_out = 8'h2F;
                    16'hD080: data_out = 8'hD0;
                    16'hD081: data_out = 8'hD1;
                    16'hD082: data_out = 8'hD2;
                    16'hD083: data_out = 8'hD3;
                    16'hD084: data_out = 8'hD4;
                    16'hD085: data_out = 8'hD5;
                    16'hD086: data_out = 8'hD6;
                    16'hD087: data_out = 8'hD7;
                    16'hD088: data_out = 8'hD8;
                    16'hD089: data_out = 8'hD9;
                    16'hD08A: data_out = 8'hDA;
                    16'hD08B: data_out = 8'hDB;
                    16'hD08C: data_out = 8'hDC;
                    16'hD08D: data_out = 8'hDD;
                    16'hD08E: data_out = 8'hDE;
                    16'hD08F: data_out = 8'hDF;
                    16'hD090: data_out = 8'hE0;
                    16'hD091: data_out = 8'hE1;
                    16'hD092: data_out = 8'hE2;
                    16'hD093: data_out = 8'hE3;
                    16'hD094: data_out = 8'hE4;
                    16'hD095: data_out = 8'hE5;
                    16'hD096: data_out = 8'hE6;
                    16'hD097: data_out = 8'hE7;
                    16'hD098: data_out = 8'hE8;
                    16'hD099: data_out = 8'hE9;
                    16'hD09A: data_out = 8'hEA;
                    16'hD09B: data_out = 8'hEB;
                    16'hD09C: data_out = 8'hEC;
                    16'hD09D: data_out = 8'hED;
                    16'hD09E: data_out = 8'hEE;
                    16'hD09F: data_out = 8'hEF;
                    16'hD0A0: data_out = 8'hF0;
                    16'hD0A1: data_out = 8'hF1;
                    16'hD0A2: data_out = 8'hF2;
                    16'hD0A3: data_out = 8'hF3;
                    16'hD0A4: data_out = 8'hF4;
                    16'hD0A5: data_out = 8'hF5;
                    16'hD0A6: data_out = 8'hF6;
                    16'hD0A7: data_out = 8'hF7;
                    16'hD0A8: data_out = 8'hF8;
                    16'hD0A9: data_out = 8'hF9;
                    16'hD0AA: data_out = 8'hFA;
                    16'hD0AB: data_out = 8'hFB;
                    16'hD0AC: data_out = 8'hFC;
                    16'hD0AD: data_out = 8'hFD;
                    16'hD0AE: data_out = 8'hFE;
                    16'hD0AF: data_out = 8'hFF;
                    16'hD0B0: data_out = 8'h80;
                    16'hD0B1: data_out = 8'h81;
                    16'hD0B2: data_out = 8'h82;
                    16'hD0B3: data_out = 8'h83;
                    16'hD0B4: data_out = 8'h84;
                    16'hD0B5: data_out = 8'h85;
                    16'hD0B6: data_out = 8'h86;
                    16'hD0B7: data_out = 8'h87;
                    16'hD0B8: data_out = 8'h88;
                    16'hD0B9: data_out = 8'h89;
                    16'hD0BA: data_out = 8'h8A;
                    16'hD0BB: data_out = 8'h8B;
                    16'hD0BC: data_out = 8'h8C;
                    16'hD0BD: data_out = 8'h8D;
                    16'hD0BE: data_out = 8'h8E;
                    16'hD0BF: data_out = 8'h8F;
                    16'hD0C0: data_out = 8'h90;
                    16'hD0C1: data_out = 8'h91;
                    16'hD0C2: data_out = 8'h92;
                    16'hD0C3: data_out = 8'h93;
                    16'hD0C4: data_out = 8'h94;
                    16'hD0C5: data_out = 8'h95;
                    16'hD0C6: data_out = 8'h96;
                    16'hD0C7: data_out = 8'h97;
                    16'hD0C8: data_out = 8'h98;
                    16'hD0C9: data_out = 8'h99;
                    16'hD0CA: data_out = 8'h9A;
                    16'hD0CB: data_out = 8'h9B;
                    16'hD0CC: data_out = 8'h9C;
                    16'hD0CD: data_out = 8'h9D;
                    16'hD0CE: data_out = 8'h9E;
                    16'hD0CF: data_out = 8'h9F;
                    16'hD0D0: data_out = 8'hA0;
                    16'hD0D1: data_out = 8'hA1;
                    16'hD0D2: data_out = 8'hA2;
                    16'hD0D3: data_out = 8'hA3;
                    16'hD0D4: data_out = 8'hA4;
                    16'hD0D5: data_out = 8'hA5;
                    16'hD0D6: data_out = 8'hA6;
                    16'hD0D7: data_out = 8'hA7;
                    16'hD0D8: data_out = 8'hA8;
                    16'hD0D9: data_out = 8'hA9;
                    16'hD0DA: data_out = 8'hAA;
                    16'hD0DB: data_out = 8'hAB;
                    16'hD0DC: data_out = 8'hAC;
                    16'hD0DD: data_out = 8'hAD;
                    16'hD0DE: data_out = 8'hAE;
                    16'hD0DF: data_out = 8'hAF;
                    16'hD0E0: data_out = 8'hB0;
                    16'hD0E1: data_out = 8'hB1;
                    16'hD0E2: data_out = 8'hB2;
                    16'hD0E3: data_out = 8'hB3;
                    16'hD0E4: data_out = 8'hB4;
                    16'hD0E5: data_out = 8'hB5;
                    16'hD0E6: data_out = 8'hB6;
                    16'hD0E7: data_out = 8'hB7;
                    16'hD0E8: data_out = 8'hB8;
                    16'hD0E9: data_out = 8'hB9;
                    16'hD0EA: data_out = 8'hBA;
                    16'hD0EB: data_out = 8'hBB;
                    16'hD0EC: data_out = 8'hBC;
                    16'hD0ED: data_out = 8'hBD;
                    16'hD0EE: data_out = 8'hBE;
                    16'hD0EF: data_out = 8'hBF;
                    16'hD0F0: data_out = 8'hC0;
                    16'hD0F1: data_out = 8'hC1;
                    16'hD0F2: data_out = 8'hC2;
                    16'hD0F3: data_out = 8'hC3;
                    16'hD0F4: data_out = 8'hC4;
                    16'hD0F5: data_out = 8'hC5;
                    16'hD0F6: data_out = 8'hC6;
                    16'hD0F7: data_out = 8'hC7;
                    16'hD0F8: data_out = 8'hC8;
                    16'hD0F9: data_out = 8'hC9;
                    16'hD0FA: data_out = 8'hCA;
                    16'hD0FB: data_out = 8'hCB;
                    16'hD0FC: data_out = 8'hCC;
                    16'hD0FD: data_out = 8'hCD;
                    16'hD0FE: data_out = 8'hCE;
                    16'hD0FF: data_out = 8'hCF;
                    16'hD100: data_out = 8'hD1;
                    16'hD101: data_out = 8'hD0;
                    16'hD102: data_out = 8'hCF;
                    16'hD103: data_out = 8'hCE;
                    16'hD104: data_out = 8'hCD;
                    16'hD105: data_out = 8'hCC;
                    16'hD106: data_out = 8'hCB;
                    16'hD107: data_out = 8'hCA;
                    16'hD108: data_out = 8'hC9;
                    16'hD109: data_out = 8'hC8;
                    16'hD10A: data_out = 8'hC7;
                    16'hD10B: data_out = 8'hC6;
                    16'hD10C: data_out = 8'hC5;
                    16'hD10D: data_out = 8'hC4;
                    16'hD10E: data_out = 8'hC3;
                    16'hD10F: data_out = 8'hC2;
                    16'hD110: data_out = 8'hC1;
                    16'hD111: data_out = 8'hC0;
                    16'hD112: data_out = 8'hBF;
                    16'hD113: data_out = 8'hBE;
                    16'hD114: data_out = 8'hBD;
                    16'hD115: data_out = 8'hBC;
                    16'hD116: data_out = 8'hBB;
                    16'hD117: data_out = 8'hBA;
                    16'hD118: data_out = 8'hB9;
                    16'hD119: data_out = 8'hB8;
                    16'hD11A: data_out = 8'hB7;
                    16'hD11B: data_out = 8'hB6;
                    16'hD11C: data_out = 8'hB5;
                    16'hD11D: data_out = 8'hB4;
                    16'hD11E: data_out = 8'hB3;
                    16'hD11F: data_out = 8'hB2;
                    16'hD120: data_out = 8'hB1;
                    16'hD121: data_out = 8'hB0;
                    16'hD122: data_out = 8'hAF;
                    16'hD123: data_out = 8'hAE;
                    16'hD124: data_out = 8'hAD;
                    16'hD125: data_out = 8'hAC;
                    16'hD126: data_out = 8'hAB;
                    16'hD127: data_out = 8'hAA;
                    16'hD128: data_out = 8'hA9;
                    16'hD129: data_out = 8'hA8;
                    16'hD12A: data_out = 8'hA7;
                    16'hD12B: data_out = 8'hA6;
                    16'hD12C: data_out = 8'hA5;
                    16'hD12D: data_out = 8'hA4;
                    16'hD12E: data_out = 8'hA3;
                    16'hD12F: data_out = 8'hA2;
                    16'hD130: data_out = 8'hA1;
                    16'hD131: data_out = 8'hA0;
                    16'hD132: data_out = 8'h9F;
                    16'hD133: data_out = 8'h9E;
                    16'hD134: data_out = 8'h9D;
                    16'hD135: data_out = 8'h9C;
                    16'hD136: data_out = 8'h9B;
                    16'hD137: data_out = 8'h9A;
                    16'hD138: data_out = 8'h99;
                    16'hD139: data_out = 8'h98;
                    16'hD13A: data_out = 8'h97;
                    16'hD13B: data_out = 8'h96;
                    16'hD13C: data_out = 8'h95;
                    16'hD13D: data_out = 8'h94;
                    16'hD13E: data_out = 8'h93;
                    16'hD13F: data_out = 8'h92;
                    16'hD140: data_out = 8'h91;
                    16'hD141: data_out = 8'h90;
                    16'hD142: data_out = 8'h8F;
                    16'hD143: data_out = 8'h8E;
                    16'hD144: data_out = 8'h8D;
                    16'hD145: data_out = 8'h8C;
                    16'hD146: data_out = 8'h8B;
                    16'hD147: data_out = 8'h8A;
                    16'hD148: data_out = 8'h89;
                    16'hD149: data_out = 8'h88;
                    16'hD14A: data_out = 8'h87;
                    16'hD14B: data_out = 8'h86;
                    16'hD14C: data_out = 8'h85;
                    16'hD14D: data_out = 8'h84;
                    16'hD14E: data_out = 8'h83;
                    16'hD14F: data_out = 8'h82;
                    16'hD150: data_out = 8'h81;
                    16'hD151: data_out = 8'h0;
                    16'hD152: data_out = 8'h1;
                    16'hD153: data_out = 8'h2;
                    16'hD154: data_out = 8'h3;
                    16'hD155: data_out = 8'h4;
                    16'hD156: data_out = 8'h5;
                    16'hD157: data_out = 8'h6;
                    16'hD158: data_out = 8'h7;
                    16'hD159: data_out = 8'h8;
                    16'hD15A: data_out = 8'h9;
                    16'hD15B: data_out = 8'hA;
                    16'hD15C: data_out = 8'hB;
                    16'hD15D: data_out = 8'hC;
                    16'hD15E: data_out = 8'hD;
                    16'hD15F: data_out = 8'hE;
                    16'hD160: data_out = 8'hF;
                    16'hD161: data_out = 8'h10;
                    16'hD162: data_out = 8'h11;
                    16'hD163: data_out = 8'h12;
                    16'hD164: data_out = 8'h13;
                    16'hD165: data_out = 8'h14;
                    16'hD166: data_out = 8'h15;
                    16'hD167: data_out = 8'h16;
                    16'hD168: data_out = 8'h17;
                    16'hD169: data_out = 8'h18;
                    16'hD16A: data_out = 8'h19;
                    16'hD16B: data_out = 8'h1A;
                    16'hD16C: data_out = 8'h1B;
                    16'hD16D: data_out = 8'h1C;
                    16'hD16E: data_out = 8'h1D;
                    16'hD16F: data_out = 8'h1E;
                    16'hD170: data_out = 8'h1F;
                    16'hD171: data_out = 8'h20;
                    16'hD172: data_out = 8'h21;
                    16'hD173: data_out = 8'h22;
                    16'hD174: data_out = 8'h23;
                    16'hD175: data_out = 8'h24;
                    16'hD176: data_out = 8'h25;
                    16'hD177: data_out = 8'h26;
                    16'hD178: data_out = 8'h27;
                    16'hD179: data_out = 8'h28;
                    16'hD17A: data_out = 8'h29;
                    16'hD17B: data_out = 8'h2A;
                    16'hD17C: data_out = 8'h2B;
                    16'hD17D: data_out = 8'h2C;
                    16'hD17E: data_out = 8'h2D;
                    16'hD17F: data_out = 8'h2E;
                    16'hD180: data_out = 8'hD1;
                    16'hD181: data_out = 8'hD2;
                    16'hD182: data_out = 8'hD3;
                    16'hD183: data_out = 8'hD4;
                    16'hD184: data_out = 8'hD5;
                    16'hD185: data_out = 8'hD6;
                    16'hD186: data_out = 8'hD7;
                    16'hD187: data_out = 8'hD8;
                    16'hD188: data_out = 8'hD9;
                    16'hD189: data_out = 8'hDA;
                    16'hD18A: data_out = 8'hDB;
                    16'hD18B: data_out = 8'hDC;
                    16'hD18C: data_out = 8'hDD;
                    16'hD18D: data_out = 8'hDE;
                    16'hD18E: data_out = 8'hDF;
                    16'hD18F: data_out = 8'hE0;
                    16'hD190: data_out = 8'hE1;
                    16'hD191: data_out = 8'hE2;
                    16'hD192: data_out = 8'hE3;
                    16'hD193: data_out = 8'hE4;
                    16'hD194: data_out = 8'hE5;
                    16'hD195: data_out = 8'hE6;
                    16'hD196: data_out = 8'hE7;
                    16'hD197: data_out = 8'hE8;
                    16'hD198: data_out = 8'hE9;
                    16'hD199: data_out = 8'hEA;
                    16'hD19A: data_out = 8'hEB;
                    16'hD19B: data_out = 8'hEC;
                    16'hD19C: data_out = 8'hED;
                    16'hD19D: data_out = 8'hEE;
                    16'hD19E: data_out = 8'hEF;
                    16'hD19F: data_out = 8'hF0;
                    16'hD1A0: data_out = 8'hF1;
                    16'hD1A1: data_out = 8'hF2;
                    16'hD1A2: data_out = 8'hF3;
                    16'hD1A3: data_out = 8'hF4;
                    16'hD1A4: data_out = 8'hF5;
                    16'hD1A5: data_out = 8'hF6;
                    16'hD1A6: data_out = 8'hF7;
                    16'hD1A7: data_out = 8'hF8;
                    16'hD1A8: data_out = 8'hF9;
                    16'hD1A9: data_out = 8'hFA;
                    16'hD1AA: data_out = 8'hFB;
                    16'hD1AB: data_out = 8'hFC;
                    16'hD1AC: data_out = 8'hFD;
                    16'hD1AD: data_out = 8'hFE;
                    16'hD1AE: data_out = 8'hFF;
                    16'hD1AF: data_out = 8'h80;
                    16'hD1B0: data_out = 8'h81;
                    16'hD1B1: data_out = 8'h82;
                    16'hD1B2: data_out = 8'h83;
                    16'hD1B3: data_out = 8'h84;
                    16'hD1B4: data_out = 8'h85;
                    16'hD1B5: data_out = 8'h86;
                    16'hD1B6: data_out = 8'h87;
                    16'hD1B7: data_out = 8'h88;
                    16'hD1B8: data_out = 8'h89;
                    16'hD1B9: data_out = 8'h8A;
                    16'hD1BA: data_out = 8'h8B;
                    16'hD1BB: data_out = 8'h8C;
                    16'hD1BC: data_out = 8'h8D;
                    16'hD1BD: data_out = 8'h8E;
                    16'hD1BE: data_out = 8'h8F;
                    16'hD1BF: data_out = 8'h90;
                    16'hD1C0: data_out = 8'h91;
                    16'hD1C1: data_out = 8'h92;
                    16'hD1C2: data_out = 8'h93;
                    16'hD1C3: data_out = 8'h94;
                    16'hD1C4: data_out = 8'h95;
                    16'hD1C5: data_out = 8'h96;
                    16'hD1C6: data_out = 8'h97;
                    16'hD1C7: data_out = 8'h98;
                    16'hD1C8: data_out = 8'h99;
                    16'hD1C9: data_out = 8'h9A;
                    16'hD1CA: data_out = 8'h9B;
                    16'hD1CB: data_out = 8'h9C;
                    16'hD1CC: data_out = 8'h9D;
                    16'hD1CD: data_out = 8'h9E;
                    16'hD1CE: data_out = 8'h9F;
                    16'hD1CF: data_out = 8'hA0;
                    16'hD1D0: data_out = 8'hA1;
                    16'hD1D1: data_out = 8'hA2;
                    16'hD1D2: data_out = 8'hA3;
                    16'hD1D3: data_out = 8'hA4;
                    16'hD1D4: data_out = 8'hA5;
                    16'hD1D5: data_out = 8'hA6;
                    16'hD1D6: data_out = 8'hA7;
                    16'hD1D7: data_out = 8'hA8;
                    16'hD1D8: data_out = 8'hA9;
                    16'hD1D9: data_out = 8'hAA;
                    16'hD1DA: data_out = 8'hAB;
                    16'hD1DB: data_out = 8'hAC;
                    16'hD1DC: data_out = 8'hAD;
                    16'hD1DD: data_out = 8'hAE;
                    16'hD1DE: data_out = 8'hAF;
                    16'hD1DF: data_out = 8'hB0;
                    16'hD1E0: data_out = 8'hB1;
                    16'hD1E1: data_out = 8'hB2;
                    16'hD1E2: data_out = 8'hB3;
                    16'hD1E3: data_out = 8'hB4;
                    16'hD1E4: data_out = 8'hB5;
                    16'hD1E5: data_out = 8'hB6;
                    16'hD1E6: data_out = 8'hB7;
                    16'hD1E7: data_out = 8'hB8;
                    16'hD1E8: data_out = 8'hB9;
                    16'hD1E9: data_out = 8'hBA;
                    16'hD1EA: data_out = 8'hBB;
                    16'hD1EB: data_out = 8'hBC;
                    16'hD1EC: data_out = 8'hBD;
                    16'hD1ED: data_out = 8'hBE;
                    16'hD1EE: data_out = 8'hBF;
                    16'hD1EF: data_out = 8'hC0;
                    16'hD1F0: data_out = 8'hC1;
                    16'hD1F1: data_out = 8'hC2;
                    16'hD1F2: data_out = 8'hC3;
                    16'hD1F3: data_out = 8'hC4;
                    16'hD1F4: data_out = 8'hC5;
                    16'hD1F5: data_out = 8'hC6;
                    16'hD1F6: data_out = 8'hC7;
                    16'hD1F7: data_out = 8'hC8;
                    16'hD1F8: data_out = 8'hC9;
                    16'hD1F9: data_out = 8'hCA;
                    16'hD1FA: data_out = 8'hCB;
                    16'hD1FB: data_out = 8'hCC;
                    16'hD1FC: data_out = 8'hCD;
                    16'hD1FD: data_out = 8'hCE;
                    16'hD1FE: data_out = 8'hCF;
                    16'hD1FF: data_out = 8'hD0;
                    16'hD200: data_out = 8'hD2;
                    16'hD201: data_out = 8'hD1;
                    16'hD202: data_out = 8'hD0;
                    16'hD203: data_out = 8'hCF;
                    16'hD204: data_out = 8'hCE;
                    16'hD205: data_out = 8'hCD;
                    16'hD206: data_out = 8'hCC;
                    16'hD207: data_out = 8'hCB;
                    16'hD208: data_out = 8'hCA;
                    16'hD209: data_out = 8'hC9;
                    16'hD20A: data_out = 8'hC8;
                    16'hD20B: data_out = 8'hC7;
                    16'hD20C: data_out = 8'hC6;
                    16'hD20D: data_out = 8'hC5;
                    16'hD20E: data_out = 8'hC4;
                    16'hD20F: data_out = 8'hC3;
                    16'hD210: data_out = 8'hC2;
                    16'hD211: data_out = 8'hC1;
                    16'hD212: data_out = 8'hC0;
                    16'hD213: data_out = 8'hBF;
                    16'hD214: data_out = 8'hBE;
                    16'hD215: data_out = 8'hBD;
                    16'hD216: data_out = 8'hBC;
                    16'hD217: data_out = 8'hBB;
                    16'hD218: data_out = 8'hBA;
                    16'hD219: data_out = 8'hB9;
                    16'hD21A: data_out = 8'hB8;
                    16'hD21B: data_out = 8'hB7;
                    16'hD21C: data_out = 8'hB6;
                    16'hD21D: data_out = 8'hB5;
                    16'hD21E: data_out = 8'hB4;
                    16'hD21F: data_out = 8'hB3;
                    16'hD220: data_out = 8'hB2;
                    16'hD221: data_out = 8'hB1;
                    16'hD222: data_out = 8'hB0;
                    16'hD223: data_out = 8'hAF;
                    16'hD224: data_out = 8'hAE;
                    16'hD225: data_out = 8'hAD;
                    16'hD226: data_out = 8'hAC;
                    16'hD227: data_out = 8'hAB;
                    16'hD228: data_out = 8'hAA;
                    16'hD229: data_out = 8'hA9;
                    16'hD22A: data_out = 8'hA8;
                    16'hD22B: data_out = 8'hA7;
                    16'hD22C: data_out = 8'hA6;
                    16'hD22D: data_out = 8'hA5;
                    16'hD22E: data_out = 8'hA4;
                    16'hD22F: data_out = 8'hA3;
                    16'hD230: data_out = 8'hA2;
                    16'hD231: data_out = 8'hA1;
                    16'hD232: data_out = 8'hA0;
                    16'hD233: data_out = 8'h9F;
                    16'hD234: data_out = 8'h9E;
                    16'hD235: data_out = 8'h9D;
                    16'hD236: data_out = 8'h9C;
                    16'hD237: data_out = 8'h9B;
                    16'hD238: data_out = 8'h9A;
                    16'hD239: data_out = 8'h99;
                    16'hD23A: data_out = 8'h98;
                    16'hD23B: data_out = 8'h97;
                    16'hD23C: data_out = 8'h96;
                    16'hD23D: data_out = 8'h95;
                    16'hD23E: data_out = 8'h94;
                    16'hD23F: data_out = 8'h93;
                    16'hD240: data_out = 8'h92;
                    16'hD241: data_out = 8'h91;
                    16'hD242: data_out = 8'h90;
                    16'hD243: data_out = 8'h8F;
                    16'hD244: data_out = 8'h8E;
                    16'hD245: data_out = 8'h8D;
                    16'hD246: data_out = 8'h8C;
                    16'hD247: data_out = 8'h8B;
                    16'hD248: data_out = 8'h8A;
                    16'hD249: data_out = 8'h89;
                    16'hD24A: data_out = 8'h88;
                    16'hD24B: data_out = 8'h87;
                    16'hD24C: data_out = 8'h86;
                    16'hD24D: data_out = 8'h85;
                    16'hD24E: data_out = 8'h84;
                    16'hD24F: data_out = 8'h83;
                    16'hD250: data_out = 8'h82;
                    16'hD251: data_out = 8'h81;
                    16'hD252: data_out = 8'h0;
                    16'hD253: data_out = 8'h1;
                    16'hD254: data_out = 8'h2;
                    16'hD255: data_out = 8'h3;
                    16'hD256: data_out = 8'h4;
                    16'hD257: data_out = 8'h5;
                    16'hD258: data_out = 8'h6;
                    16'hD259: data_out = 8'h7;
                    16'hD25A: data_out = 8'h8;
                    16'hD25B: data_out = 8'h9;
                    16'hD25C: data_out = 8'hA;
                    16'hD25D: data_out = 8'hB;
                    16'hD25E: data_out = 8'hC;
                    16'hD25F: data_out = 8'hD;
                    16'hD260: data_out = 8'hE;
                    16'hD261: data_out = 8'hF;
                    16'hD262: data_out = 8'h10;
                    16'hD263: data_out = 8'h11;
                    16'hD264: data_out = 8'h12;
                    16'hD265: data_out = 8'h13;
                    16'hD266: data_out = 8'h14;
                    16'hD267: data_out = 8'h15;
                    16'hD268: data_out = 8'h16;
                    16'hD269: data_out = 8'h17;
                    16'hD26A: data_out = 8'h18;
                    16'hD26B: data_out = 8'h19;
                    16'hD26C: data_out = 8'h1A;
                    16'hD26D: data_out = 8'h1B;
                    16'hD26E: data_out = 8'h1C;
                    16'hD26F: data_out = 8'h1D;
                    16'hD270: data_out = 8'h1E;
                    16'hD271: data_out = 8'h1F;
                    16'hD272: data_out = 8'h20;
                    16'hD273: data_out = 8'h21;
                    16'hD274: data_out = 8'h22;
                    16'hD275: data_out = 8'h23;
                    16'hD276: data_out = 8'h24;
                    16'hD277: data_out = 8'h25;
                    16'hD278: data_out = 8'h26;
                    16'hD279: data_out = 8'h27;
                    16'hD27A: data_out = 8'h28;
                    16'hD27B: data_out = 8'h29;
                    16'hD27C: data_out = 8'h2A;
                    16'hD27D: data_out = 8'h2B;
                    16'hD27E: data_out = 8'h2C;
                    16'hD27F: data_out = 8'h2D;
                    16'hD280: data_out = 8'hD2;
                    16'hD281: data_out = 8'hD3;
                    16'hD282: data_out = 8'hD4;
                    16'hD283: data_out = 8'hD5;
                    16'hD284: data_out = 8'hD6;
                    16'hD285: data_out = 8'hD7;
                    16'hD286: data_out = 8'hD8;
                    16'hD287: data_out = 8'hD9;
                    16'hD288: data_out = 8'hDA;
                    16'hD289: data_out = 8'hDB;
                    16'hD28A: data_out = 8'hDC;
                    16'hD28B: data_out = 8'hDD;
                    16'hD28C: data_out = 8'hDE;
                    16'hD28D: data_out = 8'hDF;
                    16'hD28E: data_out = 8'hE0;
                    16'hD28F: data_out = 8'hE1;
                    16'hD290: data_out = 8'hE2;
                    16'hD291: data_out = 8'hE3;
                    16'hD292: data_out = 8'hE4;
                    16'hD293: data_out = 8'hE5;
                    16'hD294: data_out = 8'hE6;
                    16'hD295: data_out = 8'hE7;
                    16'hD296: data_out = 8'hE8;
                    16'hD297: data_out = 8'hE9;
                    16'hD298: data_out = 8'hEA;
                    16'hD299: data_out = 8'hEB;
                    16'hD29A: data_out = 8'hEC;
                    16'hD29B: data_out = 8'hED;
                    16'hD29C: data_out = 8'hEE;
                    16'hD29D: data_out = 8'hEF;
                    16'hD29E: data_out = 8'hF0;
                    16'hD29F: data_out = 8'hF1;
                    16'hD2A0: data_out = 8'hF2;
                    16'hD2A1: data_out = 8'hF3;
                    16'hD2A2: data_out = 8'hF4;
                    16'hD2A3: data_out = 8'hF5;
                    16'hD2A4: data_out = 8'hF6;
                    16'hD2A5: data_out = 8'hF7;
                    16'hD2A6: data_out = 8'hF8;
                    16'hD2A7: data_out = 8'hF9;
                    16'hD2A8: data_out = 8'hFA;
                    16'hD2A9: data_out = 8'hFB;
                    16'hD2AA: data_out = 8'hFC;
                    16'hD2AB: data_out = 8'hFD;
                    16'hD2AC: data_out = 8'hFE;
                    16'hD2AD: data_out = 8'hFF;
                    16'hD2AE: data_out = 8'h80;
                    16'hD2AF: data_out = 8'h81;
                    16'hD2B0: data_out = 8'h82;
                    16'hD2B1: data_out = 8'h83;
                    16'hD2B2: data_out = 8'h84;
                    16'hD2B3: data_out = 8'h85;
                    16'hD2B4: data_out = 8'h86;
                    16'hD2B5: data_out = 8'h87;
                    16'hD2B6: data_out = 8'h88;
                    16'hD2B7: data_out = 8'h89;
                    16'hD2B8: data_out = 8'h8A;
                    16'hD2B9: data_out = 8'h8B;
                    16'hD2BA: data_out = 8'h8C;
                    16'hD2BB: data_out = 8'h8D;
                    16'hD2BC: data_out = 8'h8E;
                    16'hD2BD: data_out = 8'h8F;
                    16'hD2BE: data_out = 8'h90;
                    16'hD2BF: data_out = 8'h91;
                    16'hD2C0: data_out = 8'h92;
                    16'hD2C1: data_out = 8'h93;
                    16'hD2C2: data_out = 8'h94;
                    16'hD2C3: data_out = 8'h95;
                    16'hD2C4: data_out = 8'h96;
                    16'hD2C5: data_out = 8'h97;
                    16'hD2C6: data_out = 8'h98;
                    16'hD2C7: data_out = 8'h99;
                    16'hD2C8: data_out = 8'h9A;
                    16'hD2C9: data_out = 8'h9B;
                    16'hD2CA: data_out = 8'h9C;
                    16'hD2CB: data_out = 8'h9D;
                    16'hD2CC: data_out = 8'h9E;
                    16'hD2CD: data_out = 8'h9F;
                    16'hD2CE: data_out = 8'hA0;
                    16'hD2CF: data_out = 8'hA1;
                    16'hD2D0: data_out = 8'hA2;
                    16'hD2D1: data_out = 8'hA3;
                    16'hD2D2: data_out = 8'hA4;
                    16'hD2D3: data_out = 8'hA5;
                    16'hD2D4: data_out = 8'hA6;
                    16'hD2D5: data_out = 8'hA7;
                    16'hD2D6: data_out = 8'hA8;
                    16'hD2D7: data_out = 8'hA9;
                    16'hD2D8: data_out = 8'hAA;
                    16'hD2D9: data_out = 8'hAB;
                    16'hD2DA: data_out = 8'hAC;
                    16'hD2DB: data_out = 8'hAD;
                    16'hD2DC: data_out = 8'hAE;
                    16'hD2DD: data_out = 8'hAF;
                    16'hD2DE: data_out = 8'hB0;
                    16'hD2DF: data_out = 8'hB1;
                    16'hD2E0: data_out = 8'hB2;
                    16'hD2E1: data_out = 8'hB3;
                    16'hD2E2: data_out = 8'hB4;
                    16'hD2E3: data_out = 8'hB5;
                    16'hD2E4: data_out = 8'hB6;
                    16'hD2E5: data_out = 8'hB7;
                    16'hD2E6: data_out = 8'hB8;
                    16'hD2E7: data_out = 8'hB9;
                    16'hD2E8: data_out = 8'hBA;
                    16'hD2E9: data_out = 8'hBB;
                    16'hD2EA: data_out = 8'hBC;
                    16'hD2EB: data_out = 8'hBD;
                    16'hD2EC: data_out = 8'hBE;
                    16'hD2ED: data_out = 8'hBF;
                    16'hD2EE: data_out = 8'hC0;
                    16'hD2EF: data_out = 8'hC1;
                    16'hD2F0: data_out = 8'hC2;
                    16'hD2F1: data_out = 8'hC3;
                    16'hD2F2: data_out = 8'hC4;
                    16'hD2F3: data_out = 8'hC5;
                    16'hD2F4: data_out = 8'hC6;
                    16'hD2F5: data_out = 8'hC7;
                    16'hD2F6: data_out = 8'hC8;
                    16'hD2F7: data_out = 8'hC9;
                    16'hD2F8: data_out = 8'hCA;
                    16'hD2F9: data_out = 8'hCB;
                    16'hD2FA: data_out = 8'hCC;
                    16'hD2FB: data_out = 8'hCD;
                    16'hD2FC: data_out = 8'hCE;
                    16'hD2FD: data_out = 8'hCF;
                    16'hD2FE: data_out = 8'hD0;
                    16'hD2FF: data_out = 8'hD1;
                    16'hD300: data_out = 8'hD3;
                    16'hD301: data_out = 8'hD2;
                    16'hD302: data_out = 8'hD1;
                    16'hD303: data_out = 8'hD0;
                    16'hD304: data_out = 8'hCF;
                    16'hD305: data_out = 8'hCE;
                    16'hD306: data_out = 8'hCD;
                    16'hD307: data_out = 8'hCC;
                    16'hD308: data_out = 8'hCB;
                    16'hD309: data_out = 8'hCA;
                    16'hD30A: data_out = 8'hC9;
                    16'hD30B: data_out = 8'hC8;
                    16'hD30C: data_out = 8'hC7;
                    16'hD30D: data_out = 8'hC6;
                    16'hD30E: data_out = 8'hC5;
                    16'hD30F: data_out = 8'hC4;
                    16'hD310: data_out = 8'hC3;
                    16'hD311: data_out = 8'hC2;
                    16'hD312: data_out = 8'hC1;
                    16'hD313: data_out = 8'hC0;
                    16'hD314: data_out = 8'hBF;
                    16'hD315: data_out = 8'hBE;
                    16'hD316: data_out = 8'hBD;
                    16'hD317: data_out = 8'hBC;
                    16'hD318: data_out = 8'hBB;
                    16'hD319: data_out = 8'hBA;
                    16'hD31A: data_out = 8'hB9;
                    16'hD31B: data_out = 8'hB8;
                    16'hD31C: data_out = 8'hB7;
                    16'hD31D: data_out = 8'hB6;
                    16'hD31E: data_out = 8'hB5;
                    16'hD31F: data_out = 8'hB4;
                    16'hD320: data_out = 8'hB3;
                    16'hD321: data_out = 8'hB2;
                    16'hD322: data_out = 8'hB1;
                    16'hD323: data_out = 8'hB0;
                    16'hD324: data_out = 8'hAF;
                    16'hD325: data_out = 8'hAE;
                    16'hD326: data_out = 8'hAD;
                    16'hD327: data_out = 8'hAC;
                    16'hD328: data_out = 8'hAB;
                    16'hD329: data_out = 8'hAA;
                    16'hD32A: data_out = 8'hA9;
                    16'hD32B: data_out = 8'hA8;
                    16'hD32C: data_out = 8'hA7;
                    16'hD32D: data_out = 8'hA6;
                    16'hD32E: data_out = 8'hA5;
                    16'hD32F: data_out = 8'hA4;
                    16'hD330: data_out = 8'hA3;
                    16'hD331: data_out = 8'hA2;
                    16'hD332: data_out = 8'hA1;
                    16'hD333: data_out = 8'hA0;
                    16'hD334: data_out = 8'h9F;
                    16'hD335: data_out = 8'h9E;
                    16'hD336: data_out = 8'h9D;
                    16'hD337: data_out = 8'h9C;
                    16'hD338: data_out = 8'h9B;
                    16'hD339: data_out = 8'h9A;
                    16'hD33A: data_out = 8'h99;
                    16'hD33B: data_out = 8'h98;
                    16'hD33C: data_out = 8'h97;
                    16'hD33D: data_out = 8'h96;
                    16'hD33E: data_out = 8'h95;
                    16'hD33F: data_out = 8'h94;
                    16'hD340: data_out = 8'h93;
                    16'hD341: data_out = 8'h92;
                    16'hD342: data_out = 8'h91;
                    16'hD343: data_out = 8'h90;
                    16'hD344: data_out = 8'h8F;
                    16'hD345: data_out = 8'h8E;
                    16'hD346: data_out = 8'h8D;
                    16'hD347: data_out = 8'h8C;
                    16'hD348: data_out = 8'h8B;
                    16'hD349: data_out = 8'h8A;
                    16'hD34A: data_out = 8'h89;
                    16'hD34B: data_out = 8'h88;
                    16'hD34C: data_out = 8'h87;
                    16'hD34D: data_out = 8'h86;
                    16'hD34E: data_out = 8'h85;
                    16'hD34F: data_out = 8'h84;
                    16'hD350: data_out = 8'h83;
                    16'hD351: data_out = 8'h82;
                    16'hD352: data_out = 8'h81;
                    16'hD353: data_out = 8'h0;
                    16'hD354: data_out = 8'h1;
                    16'hD355: data_out = 8'h2;
                    16'hD356: data_out = 8'h3;
                    16'hD357: data_out = 8'h4;
                    16'hD358: data_out = 8'h5;
                    16'hD359: data_out = 8'h6;
                    16'hD35A: data_out = 8'h7;
                    16'hD35B: data_out = 8'h8;
                    16'hD35C: data_out = 8'h9;
                    16'hD35D: data_out = 8'hA;
                    16'hD35E: data_out = 8'hB;
                    16'hD35F: data_out = 8'hC;
                    16'hD360: data_out = 8'hD;
                    16'hD361: data_out = 8'hE;
                    16'hD362: data_out = 8'hF;
                    16'hD363: data_out = 8'h10;
                    16'hD364: data_out = 8'h11;
                    16'hD365: data_out = 8'h12;
                    16'hD366: data_out = 8'h13;
                    16'hD367: data_out = 8'h14;
                    16'hD368: data_out = 8'h15;
                    16'hD369: data_out = 8'h16;
                    16'hD36A: data_out = 8'h17;
                    16'hD36B: data_out = 8'h18;
                    16'hD36C: data_out = 8'h19;
                    16'hD36D: data_out = 8'h1A;
                    16'hD36E: data_out = 8'h1B;
                    16'hD36F: data_out = 8'h1C;
                    16'hD370: data_out = 8'h1D;
                    16'hD371: data_out = 8'h1E;
                    16'hD372: data_out = 8'h1F;
                    16'hD373: data_out = 8'h20;
                    16'hD374: data_out = 8'h21;
                    16'hD375: data_out = 8'h22;
                    16'hD376: data_out = 8'h23;
                    16'hD377: data_out = 8'h24;
                    16'hD378: data_out = 8'h25;
                    16'hD379: data_out = 8'h26;
                    16'hD37A: data_out = 8'h27;
                    16'hD37B: data_out = 8'h28;
                    16'hD37C: data_out = 8'h29;
                    16'hD37D: data_out = 8'h2A;
                    16'hD37E: data_out = 8'h2B;
                    16'hD37F: data_out = 8'h2C;
                    16'hD380: data_out = 8'hD3;
                    16'hD381: data_out = 8'hD4;
                    16'hD382: data_out = 8'hD5;
                    16'hD383: data_out = 8'hD6;
                    16'hD384: data_out = 8'hD7;
                    16'hD385: data_out = 8'hD8;
                    16'hD386: data_out = 8'hD9;
                    16'hD387: data_out = 8'hDA;
                    16'hD388: data_out = 8'hDB;
                    16'hD389: data_out = 8'hDC;
                    16'hD38A: data_out = 8'hDD;
                    16'hD38B: data_out = 8'hDE;
                    16'hD38C: data_out = 8'hDF;
                    16'hD38D: data_out = 8'hE0;
                    16'hD38E: data_out = 8'hE1;
                    16'hD38F: data_out = 8'hE2;
                    16'hD390: data_out = 8'hE3;
                    16'hD391: data_out = 8'hE4;
                    16'hD392: data_out = 8'hE5;
                    16'hD393: data_out = 8'hE6;
                    16'hD394: data_out = 8'hE7;
                    16'hD395: data_out = 8'hE8;
                    16'hD396: data_out = 8'hE9;
                    16'hD397: data_out = 8'hEA;
                    16'hD398: data_out = 8'hEB;
                    16'hD399: data_out = 8'hEC;
                    16'hD39A: data_out = 8'hED;
                    16'hD39B: data_out = 8'hEE;
                    16'hD39C: data_out = 8'hEF;
                    16'hD39D: data_out = 8'hF0;
                    16'hD39E: data_out = 8'hF1;
                    16'hD39F: data_out = 8'hF2;
                    16'hD3A0: data_out = 8'hF3;
                    16'hD3A1: data_out = 8'hF4;
                    16'hD3A2: data_out = 8'hF5;
                    16'hD3A3: data_out = 8'hF6;
                    16'hD3A4: data_out = 8'hF7;
                    16'hD3A5: data_out = 8'hF8;
                    16'hD3A6: data_out = 8'hF9;
                    16'hD3A7: data_out = 8'hFA;
                    16'hD3A8: data_out = 8'hFB;
                    16'hD3A9: data_out = 8'hFC;
                    16'hD3AA: data_out = 8'hFD;
                    16'hD3AB: data_out = 8'hFE;
                    16'hD3AC: data_out = 8'hFF;
                    16'hD3AD: data_out = 8'h80;
                    16'hD3AE: data_out = 8'h81;
                    16'hD3AF: data_out = 8'h82;
                    16'hD3B0: data_out = 8'h83;
                    16'hD3B1: data_out = 8'h84;
                    16'hD3B2: data_out = 8'h85;
                    16'hD3B3: data_out = 8'h86;
                    16'hD3B4: data_out = 8'h87;
                    16'hD3B5: data_out = 8'h88;
                    16'hD3B6: data_out = 8'h89;
                    16'hD3B7: data_out = 8'h8A;
                    16'hD3B8: data_out = 8'h8B;
                    16'hD3B9: data_out = 8'h8C;
                    16'hD3BA: data_out = 8'h8D;
                    16'hD3BB: data_out = 8'h8E;
                    16'hD3BC: data_out = 8'h8F;
                    16'hD3BD: data_out = 8'h90;
                    16'hD3BE: data_out = 8'h91;
                    16'hD3BF: data_out = 8'h92;
                    16'hD3C0: data_out = 8'h93;
                    16'hD3C1: data_out = 8'h94;
                    16'hD3C2: data_out = 8'h95;
                    16'hD3C3: data_out = 8'h96;
                    16'hD3C4: data_out = 8'h97;
                    16'hD3C5: data_out = 8'h98;
                    16'hD3C6: data_out = 8'h99;
                    16'hD3C7: data_out = 8'h9A;
                    16'hD3C8: data_out = 8'h9B;
                    16'hD3C9: data_out = 8'h9C;
                    16'hD3CA: data_out = 8'h9D;
                    16'hD3CB: data_out = 8'h9E;
                    16'hD3CC: data_out = 8'h9F;
                    16'hD3CD: data_out = 8'hA0;
                    16'hD3CE: data_out = 8'hA1;
                    16'hD3CF: data_out = 8'hA2;
                    16'hD3D0: data_out = 8'hA3;
                    16'hD3D1: data_out = 8'hA4;
                    16'hD3D2: data_out = 8'hA5;
                    16'hD3D3: data_out = 8'hA6;
                    16'hD3D4: data_out = 8'hA7;
                    16'hD3D5: data_out = 8'hA8;
                    16'hD3D6: data_out = 8'hA9;
                    16'hD3D7: data_out = 8'hAA;
                    16'hD3D8: data_out = 8'hAB;
                    16'hD3D9: data_out = 8'hAC;
                    16'hD3DA: data_out = 8'hAD;
                    16'hD3DB: data_out = 8'hAE;
                    16'hD3DC: data_out = 8'hAF;
                    16'hD3DD: data_out = 8'hB0;
                    16'hD3DE: data_out = 8'hB1;
                    16'hD3DF: data_out = 8'hB2;
                    16'hD3E0: data_out = 8'hB3;
                    16'hD3E1: data_out = 8'hB4;
                    16'hD3E2: data_out = 8'hB5;
                    16'hD3E3: data_out = 8'hB6;
                    16'hD3E4: data_out = 8'hB7;
                    16'hD3E5: data_out = 8'hB8;
                    16'hD3E6: data_out = 8'hB9;
                    16'hD3E7: data_out = 8'hBA;
                    16'hD3E8: data_out = 8'hBB;
                    16'hD3E9: data_out = 8'hBC;
                    16'hD3EA: data_out = 8'hBD;
                    16'hD3EB: data_out = 8'hBE;
                    16'hD3EC: data_out = 8'hBF;
                    16'hD3ED: data_out = 8'hC0;
                    16'hD3EE: data_out = 8'hC1;
                    16'hD3EF: data_out = 8'hC2;
                    16'hD3F0: data_out = 8'hC3;
                    16'hD3F1: data_out = 8'hC4;
                    16'hD3F2: data_out = 8'hC5;
                    16'hD3F3: data_out = 8'hC6;
                    16'hD3F4: data_out = 8'hC7;
                    16'hD3F5: data_out = 8'hC8;
                    16'hD3F6: data_out = 8'hC9;
                    16'hD3F7: data_out = 8'hCA;
                    16'hD3F8: data_out = 8'hCB;
                    16'hD3F9: data_out = 8'hCC;
                    16'hD3FA: data_out = 8'hCD;
                    16'hD3FB: data_out = 8'hCE;
                    16'hD3FC: data_out = 8'hCF;
                    16'hD3FD: data_out = 8'hD0;
                    16'hD3FE: data_out = 8'hD1;
                    16'hD3FF: data_out = 8'hD2;
                    16'hD400: data_out = 8'hD4;
                    16'hD401: data_out = 8'hD3;
                    16'hD402: data_out = 8'hD2;
                    16'hD403: data_out = 8'hD1;
                    16'hD404: data_out = 8'hD0;
                    16'hD405: data_out = 8'hCF;
                    16'hD406: data_out = 8'hCE;
                    16'hD407: data_out = 8'hCD;
                    16'hD408: data_out = 8'hCC;
                    16'hD409: data_out = 8'hCB;
                    16'hD40A: data_out = 8'hCA;
                    16'hD40B: data_out = 8'hC9;
                    16'hD40C: data_out = 8'hC8;
                    16'hD40D: data_out = 8'hC7;
                    16'hD40E: data_out = 8'hC6;
                    16'hD40F: data_out = 8'hC5;
                    16'hD410: data_out = 8'hC4;
                    16'hD411: data_out = 8'hC3;
                    16'hD412: data_out = 8'hC2;
                    16'hD413: data_out = 8'hC1;
                    16'hD414: data_out = 8'hC0;
                    16'hD415: data_out = 8'hBF;
                    16'hD416: data_out = 8'hBE;
                    16'hD417: data_out = 8'hBD;
                    16'hD418: data_out = 8'hBC;
                    16'hD419: data_out = 8'hBB;
                    16'hD41A: data_out = 8'hBA;
                    16'hD41B: data_out = 8'hB9;
                    16'hD41C: data_out = 8'hB8;
                    16'hD41D: data_out = 8'hB7;
                    16'hD41E: data_out = 8'hB6;
                    16'hD41F: data_out = 8'hB5;
                    16'hD420: data_out = 8'hB4;
                    16'hD421: data_out = 8'hB3;
                    16'hD422: data_out = 8'hB2;
                    16'hD423: data_out = 8'hB1;
                    16'hD424: data_out = 8'hB0;
                    16'hD425: data_out = 8'hAF;
                    16'hD426: data_out = 8'hAE;
                    16'hD427: data_out = 8'hAD;
                    16'hD428: data_out = 8'hAC;
                    16'hD429: data_out = 8'hAB;
                    16'hD42A: data_out = 8'hAA;
                    16'hD42B: data_out = 8'hA9;
                    16'hD42C: data_out = 8'hA8;
                    16'hD42D: data_out = 8'hA7;
                    16'hD42E: data_out = 8'hA6;
                    16'hD42F: data_out = 8'hA5;
                    16'hD430: data_out = 8'hA4;
                    16'hD431: data_out = 8'hA3;
                    16'hD432: data_out = 8'hA2;
                    16'hD433: data_out = 8'hA1;
                    16'hD434: data_out = 8'hA0;
                    16'hD435: data_out = 8'h9F;
                    16'hD436: data_out = 8'h9E;
                    16'hD437: data_out = 8'h9D;
                    16'hD438: data_out = 8'h9C;
                    16'hD439: data_out = 8'h9B;
                    16'hD43A: data_out = 8'h9A;
                    16'hD43B: data_out = 8'h99;
                    16'hD43C: data_out = 8'h98;
                    16'hD43D: data_out = 8'h97;
                    16'hD43E: data_out = 8'h96;
                    16'hD43F: data_out = 8'h95;
                    16'hD440: data_out = 8'h94;
                    16'hD441: data_out = 8'h93;
                    16'hD442: data_out = 8'h92;
                    16'hD443: data_out = 8'h91;
                    16'hD444: data_out = 8'h90;
                    16'hD445: data_out = 8'h8F;
                    16'hD446: data_out = 8'h8E;
                    16'hD447: data_out = 8'h8D;
                    16'hD448: data_out = 8'h8C;
                    16'hD449: data_out = 8'h8B;
                    16'hD44A: data_out = 8'h8A;
                    16'hD44B: data_out = 8'h89;
                    16'hD44C: data_out = 8'h88;
                    16'hD44D: data_out = 8'h87;
                    16'hD44E: data_out = 8'h86;
                    16'hD44F: data_out = 8'h85;
                    16'hD450: data_out = 8'h84;
                    16'hD451: data_out = 8'h83;
                    16'hD452: data_out = 8'h82;
                    16'hD453: data_out = 8'h81;
                    16'hD454: data_out = 8'h0;
                    16'hD455: data_out = 8'h1;
                    16'hD456: data_out = 8'h2;
                    16'hD457: data_out = 8'h3;
                    16'hD458: data_out = 8'h4;
                    16'hD459: data_out = 8'h5;
                    16'hD45A: data_out = 8'h6;
                    16'hD45B: data_out = 8'h7;
                    16'hD45C: data_out = 8'h8;
                    16'hD45D: data_out = 8'h9;
                    16'hD45E: data_out = 8'hA;
                    16'hD45F: data_out = 8'hB;
                    16'hD460: data_out = 8'hC;
                    16'hD461: data_out = 8'hD;
                    16'hD462: data_out = 8'hE;
                    16'hD463: data_out = 8'hF;
                    16'hD464: data_out = 8'h10;
                    16'hD465: data_out = 8'h11;
                    16'hD466: data_out = 8'h12;
                    16'hD467: data_out = 8'h13;
                    16'hD468: data_out = 8'h14;
                    16'hD469: data_out = 8'h15;
                    16'hD46A: data_out = 8'h16;
                    16'hD46B: data_out = 8'h17;
                    16'hD46C: data_out = 8'h18;
                    16'hD46D: data_out = 8'h19;
                    16'hD46E: data_out = 8'h1A;
                    16'hD46F: data_out = 8'h1B;
                    16'hD470: data_out = 8'h1C;
                    16'hD471: data_out = 8'h1D;
                    16'hD472: data_out = 8'h1E;
                    16'hD473: data_out = 8'h1F;
                    16'hD474: data_out = 8'h20;
                    16'hD475: data_out = 8'h21;
                    16'hD476: data_out = 8'h22;
                    16'hD477: data_out = 8'h23;
                    16'hD478: data_out = 8'h24;
                    16'hD479: data_out = 8'h25;
                    16'hD47A: data_out = 8'h26;
                    16'hD47B: data_out = 8'h27;
                    16'hD47C: data_out = 8'h28;
                    16'hD47D: data_out = 8'h29;
                    16'hD47E: data_out = 8'h2A;
                    16'hD47F: data_out = 8'h2B;
                    16'hD480: data_out = 8'hD4;
                    16'hD481: data_out = 8'hD5;
                    16'hD482: data_out = 8'hD6;
                    16'hD483: data_out = 8'hD7;
                    16'hD484: data_out = 8'hD8;
                    16'hD485: data_out = 8'hD9;
                    16'hD486: data_out = 8'hDA;
                    16'hD487: data_out = 8'hDB;
                    16'hD488: data_out = 8'hDC;
                    16'hD489: data_out = 8'hDD;
                    16'hD48A: data_out = 8'hDE;
                    16'hD48B: data_out = 8'hDF;
                    16'hD48C: data_out = 8'hE0;
                    16'hD48D: data_out = 8'hE1;
                    16'hD48E: data_out = 8'hE2;
                    16'hD48F: data_out = 8'hE3;
                    16'hD490: data_out = 8'hE4;
                    16'hD491: data_out = 8'hE5;
                    16'hD492: data_out = 8'hE6;
                    16'hD493: data_out = 8'hE7;
                    16'hD494: data_out = 8'hE8;
                    16'hD495: data_out = 8'hE9;
                    16'hD496: data_out = 8'hEA;
                    16'hD497: data_out = 8'hEB;
                    16'hD498: data_out = 8'hEC;
                    16'hD499: data_out = 8'hED;
                    16'hD49A: data_out = 8'hEE;
                    16'hD49B: data_out = 8'hEF;
                    16'hD49C: data_out = 8'hF0;
                    16'hD49D: data_out = 8'hF1;
                    16'hD49E: data_out = 8'hF2;
                    16'hD49F: data_out = 8'hF3;
                    16'hD4A0: data_out = 8'hF4;
                    16'hD4A1: data_out = 8'hF5;
                    16'hD4A2: data_out = 8'hF6;
                    16'hD4A3: data_out = 8'hF7;
                    16'hD4A4: data_out = 8'hF8;
                    16'hD4A5: data_out = 8'hF9;
                    16'hD4A6: data_out = 8'hFA;
                    16'hD4A7: data_out = 8'hFB;
                    16'hD4A8: data_out = 8'hFC;
                    16'hD4A9: data_out = 8'hFD;
                    16'hD4AA: data_out = 8'hFE;
                    16'hD4AB: data_out = 8'hFF;
                    16'hD4AC: data_out = 8'h80;
                    16'hD4AD: data_out = 8'h81;
                    16'hD4AE: data_out = 8'h82;
                    16'hD4AF: data_out = 8'h83;
                    16'hD4B0: data_out = 8'h84;
                    16'hD4B1: data_out = 8'h85;
                    16'hD4B2: data_out = 8'h86;
                    16'hD4B3: data_out = 8'h87;
                    16'hD4B4: data_out = 8'h88;
                    16'hD4B5: data_out = 8'h89;
                    16'hD4B6: data_out = 8'h8A;
                    16'hD4B7: data_out = 8'h8B;
                    16'hD4B8: data_out = 8'h8C;
                    16'hD4B9: data_out = 8'h8D;
                    16'hD4BA: data_out = 8'h8E;
                    16'hD4BB: data_out = 8'h8F;
                    16'hD4BC: data_out = 8'h90;
                    16'hD4BD: data_out = 8'h91;
                    16'hD4BE: data_out = 8'h92;
                    16'hD4BF: data_out = 8'h93;
                    16'hD4C0: data_out = 8'h94;
                    16'hD4C1: data_out = 8'h95;
                    16'hD4C2: data_out = 8'h96;
                    16'hD4C3: data_out = 8'h97;
                    16'hD4C4: data_out = 8'h98;
                    16'hD4C5: data_out = 8'h99;
                    16'hD4C6: data_out = 8'h9A;
                    16'hD4C7: data_out = 8'h9B;
                    16'hD4C8: data_out = 8'h9C;
                    16'hD4C9: data_out = 8'h9D;
                    16'hD4CA: data_out = 8'h9E;
                    16'hD4CB: data_out = 8'h9F;
                    16'hD4CC: data_out = 8'hA0;
                    16'hD4CD: data_out = 8'hA1;
                    16'hD4CE: data_out = 8'hA2;
                    16'hD4CF: data_out = 8'hA3;
                    16'hD4D0: data_out = 8'hA4;
                    16'hD4D1: data_out = 8'hA5;
                    16'hD4D2: data_out = 8'hA6;
                    16'hD4D3: data_out = 8'hA7;
                    16'hD4D4: data_out = 8'hA8;
                    16'hD4D5: data_out = 8'hA9;
                    16'hD4D6: data_out = 8'hAA;
                    16'hD4D7: data_out = 8'hAB;
                    16'hD4D8: data_out = 8'hAC;
                    16'hD4D9: data_out = 8'hAD;
                    16'hD4DA: data_out = 8'hAE;
                    16'hD4DB: data_out = 8'hAF;
                    16'hD4DC: data_out = 8'hB0;
                    16'hD4DD: data_out = 8'hB1;
                    16'hD4DE: data_out = 8'hB2;
                    16'hD4DF: data_out = 8'hB3;
                    16'hD4E0: data_out = 8'hB4;
                    16'hD4E1: data_out = 8'hB5;
                    16'hD4E2: data_out = 8'hB6;
                    16'hD4E3: data_out = 8'hB7;
                    16'hD4E4: data_out = 8'hB8;
                    16'hD4E5: data_out = 8'hB9;
                    16'hD4E6: data_out = 8'hBA;
                    16'hD4E7: data_out = 8'hBB;
                    16'hD4E8: data_out = 8'hBC;
                    16'hD4E9: data_out = 8'hBD;
                    16'hD4EA: data_out = 8'hBE;
                    16'hD4EB: data_out = 8'hBF;
                    16'hD4EC: data_out = 8'hC0;
                    16'hD4ED: data_out = 8'hC1;
                    16'hD4EE: data_out = 8'hC2;
                    16'hD4EF: data_out = 8'hC3;
                    16'hD4F0: data_out = 8'hC4;
                    16'hD4F1: data_out = 8'hC5;
                    16'hD4F2: data_out = 8'hC6;
                    16'hD4F3: data_out = 8'hC7;
                    16'hD4F4: data_out = 8'hC8;
                    16'hD4F5: data_out = 8'hC9;
                    16'hD4F6: data_out = 8'hCA;
                    16'hD4F7: data_out = 8'hCB;
                    16'hD4F8: data_out = 8'hCC;
                    16'hD4F9: data_out = 8'hCD;
                    16'hD4FA: data_out = 8'hCE;
                    16'hD4FB: data_out = 8'hCF;
                    16'hD4FC: data_out = 8'hD0;
                    16'hD4FD: data_out = 8'hD1;
                    16'hD4FE: data_out = 8'hD2;
                    16'hD4FF: data_out = 8'hD3;
                    16'hD500: data_out = 8'hD5;
                    16'hD501: data_out = 8'hD4;
                    16'hD502: data_out = 8'hD3;
                    16'hD503: data_out = 8'hD2;
                    16'hD504: data_out = 8'hD1;
                    16'hD505: data_out = 8'hD0;
                    16'hD506: data_out = 8'hCF;
                    16'hD507: data_out = 8'hCE;
                    16'hD508: data_out = 8'hCD;
                    16'hD509: data_out = 8'hCC;
                    16'hD50A: data_out = 8'hCB;
                    16'hD50B: data_out = 8'hCA;
                    16'hD50C: data_out = 8'hC9;
                    16'hD50D: data_out = 8'hC8;
                    16'hD50E: data_out = 8'hC7;
                    16'hD50F: data_out = 8'hC6;
                    16'hD510: data_out = 8'hC5;
                    16'hD511: data_out = 8'hC4;
                    16'hD512: data_out = 8'hC3;
                    16'hD513: data_out = 8'hC2;
                    16'hD514: data_out = 8'hC1;
                    16'hD515: data_out = 8'hC0;
                    16'hD516: data_out = 8'hBF;
                    16'hD517: data_out = 8'hBE;
                    16'hD518: data_out = 8'hBD;
                    16'hD519: data_out = 8'hBC;
                    16'hD51A: data_out = 8'hBB;
                    16'hD51B: data_out = 8'hBA;
                    16'hD51C: data_out = 8'hB9;
                    16'hD51D: data_out = 8'hB8;
                    16'hD51E: data_out = 8'hB7;
                    16'hD51F: data_out = 8'hB6;
                    16'hD520: data_out = 8'hB5;
                    16'hD521: data_out = 8'hB4;
                    16'hD522: data_out = 8'hB3;
                    16'hD523: data_out = 8'hB2;
                    16'hD524: data_out = 8'hB1;
                    16'hD525: data_out = 8'hB0;
                    16'hD526: data_out = 8'hAF;
                    16'hD527: data_out = 8'hAE;
                    16'hD528: data_out = 8'hAD;
                    16'hD529: data_out = 8'hAC;
                    16'hD52A: data_out = 8'hAB;
                    16'hD52B: data_out = 8'hAA;
                    16'hD52C: data_out = 8'hA9;
                    16'hD52D: data_out = 8'hA8;
                    16'hD52E: data_out = 8'hA7;
                    16'hD52F: data_out = 8'hA6;
                    16'hD530: data_out = 8'hA5;
                    16'hD531: data_out = 8'hA4;
                    16'hD532: data_out = 8'hA3;
                    16'hD533: data_out = 8'hA2;
                    16'hD534: data_out = 8'hA1;
                    16'hD535: data_out = 8'hA0;
                    16'hD536: data_out = 8'h9F;
                    16'hD537: data_out = 8'h9E;
                    16'hD538: data_out = 8'h9D;
                    16'hD539: data_out = 8'h9C;
                    16'hD53A: data_out = 8'h9B;
                    16'hD53B: data_out = 8'h9A;
                    16'hD53C: data_out = 8'h99;
                    16'hD53D: data_out = 8'h98;
                    16'hD53E: data_out = 8'h97;
                    16'hD53F: data_out = 8'h96;
                    16'hD540: data_out = 8'h95;
                    16'hD541: data_out = 8'h94;
                    16'hD542: data_out = 8'h93;
                    16'hD543: data_out = 8'h92;
                    16'hD544: data_out = 8'h91;
                    16'hD545: data_out = 8'h90;
                    16'hD546: data_out = 8'h8F;
                    16'hD547: data_out = 8'h8E;
                    16'hD548: data_out = 8'h8D;
                    16'hD549: data_out = 8'h8C;
                    16'hD54A: data_out = 8'h8B;
                    16'hD54B: data_out = 8'h8A;
                    16'hD54C: data_out = 8'h89;
                    16'hD54D: data_out = 8'h88;
                    16'hD54E: data_out = 8'h87;
                    16'hD54F: data_out = 8'h86;
                    16'hD550: data_out = 8'h85;
                    16'hD551: data_out = 8'h84;
                    16'hD552: data_out = 8'h83;
                    16'hD553: data_out = 8'h82;
                    16'hD554: data_out = 8'h81;
                    16'hD555: data_out = 8'h0;
                    16'hD556: data_out = 8'h1;
                    16'hD557: data_out = 8'h2;
                    16'hD558: data_out = 8'h3;
                    16'hD559: data_out = 8'h4;
                    16'hD55A: data_out = 8'h5;
                    16'hD55B: data_out = 8'h6;
                    16'hD55C: data_out = 8'h7;
                    16'hD55D: data_out = 8'h8;
                    16'hD55E: data_out = 8'h9;
                    16'hD55F: data_out = 8'hA;
                    16'hD560: data_out = 8'hB;
                    16'hD561: data_out = 8'hC;
                    16'hD562: data_out = 8'hD;
                    16'hD563: data_out = 8'hE;
                    16'hD564: data_out = 8'hF;
                    16'hD565: data_out = 8'h10;
                    16'hD566: data_out = 8'h11;
                    16'hD567: data_out = 8'h12;
                    16'hD568: data_out = 8'h13;
                    16'hD569: data_out = 8'h14;
                    16'hD56A: data_out = 8'h15;
                    16'hD56B: data_out = 8'h16;
                    16'hD56C: data_out = 8'h17;
                    16'hD56D: data_out = 8'h18;
                    16'hD56E: data_out = 8'h19;
                    16'hD56F: data_out = 8'h1A;
                    16'hD570: data_out = 8'h1B;
                    16'hD571: data_out = 8'h1C;
                    16'hD572: data_out = 8'h1D;
                    16'hD573: data_out = 8'h1E;
                    16'hD574: data_out = 8'h1F;
                    16'hD575: data_out = 8'h20;
                    16'hD576: data_out = 8'h21;
                    16'hD577: data_out = 8'h22;
                    16'hD578: data_out = 8'h23;
                    16'hD579: data_out = 8'h24;
                    16'hD57A: data_out = 8'h25;
                    16'hD57B: data_out = 8'h26;
                    16'hD57C: data_out = 8'h27;
                    16'hD57D: data_out = 8'h28;
                    16'hD57E: data_out = 8'h29;
                    16'hD57F: data_out = 8'h2A;
                    16'hD580: data_out = 8'hD5;
                    16'hD581: data_out = 8'hD6;
                    16'hD582: data_out = 8'hD7;
                    16'hD583: data_out = 8'hD8;
                    16'hD584: data_out = 8'hD9;
                    16'hD585: data_out = 8'hDA;
                    16'hD586: data_out = 8'hDB;
                    16'hD587: data_out = 8'hDC;
                    16'hD588: data_out = 8'hDD;
                    16'hD589: data_out = 8'hDE;
                    16'hD58A: data_out = 8'hDF;
                    16'hD58B: data_out = 8'hE0;
                    16'hD58C: data_out = 8'hE1;
                    16'hD58D: data_out = 8'hE2;
                    16'hD58E: data_out = 8'hE3;
                    16'hD58F: data_out = 8'hE4;
                    16'hD590: data_out = 8'hE5;
                    16'hD591: data_out = 8'hE6;
                    16'hD592: data_out = 8'hE7;
                    16'hD593: data_out = 8'hE8;
                    16'hD594: data_out = 8'hE9;
                    16'hD595: data_out = 8'hEA;
                    16'hD596: data_out = 8'hEB;
                    16'hD597: data_out = 8'hEC;
                    16'hD598: data_out = 8'hED;
                    16'hD599: data_out = 8'hEE;
                    16'hD59A: data_out = 8'hEF;
                    16'hD59B: data_out = 8'hF0;
                    16'hD59C: data_out = 8'hF1;
                    16'hD59D: data_out = 8'hF2;
                    16'hD59E: data_out = 8'hF3;
                    16'hD59F: data_out = 8'hF4;
                    16'hD5A0: data_out = 8'hF5;
                    16'hD5A1: data_out = 8'hF6;
                    16'hD5A2: data_out = 8'hF7;
                    16'hD5A3: data_out = 8'hF8;
                    16'hD5A4: data_out = 8'hF9;
                    16'hD5A5: data_out = 8'hFA;
                    16'hD5A6: data_out = 8'hFB;
                    16'hD5A7: data_out = 8'hFC;
                    16'hD5A8: data_out = 8'hFD;
                    16'hD5A9: data_out = 8'hFE;
                    16'hD5AA: data_out = 8'hFF;
                    16'hD5AB: data_out = 8'h80;
                    16'hD5AC: data_out = 8'h81;
                    16'hD5AD: data_out = 8'h82;
                    16'hD5AE: data_out = 8'h83;
                    16'hD5AF: data_out = 8'h84;
                    16'hD5B0: data_out = 8'h85;
                    16'hD5B1: data_out = 8'h86;
                    16'hD5B2: data_out = 8'h87;
                    16'hD5B3: data_out = 8'h88;
                    16'hD5B4: data_out = 8'h89;
                    16'hD5B5: data_out = 8'h8A;
                    16'hD5B6: data_out = 8'h8B;
                    16'hD5B7: data_out = 8'h8C;
                    16'hD5B8: data_out = 8'h8D;
                    16'hD5B9: data_out = 8'h8E;
                    16'hD5BA: data_out = 8'h8F;
                    16'hD5BB: data_out = 8'h90;
                    16'hD5BC: data_out = 8'h91;
                    16'hD5BD: data_out = 8'h92;
                    16'hD5BE: data_out = 8'h93;
                    16'hD5BF: data_out = 8'h94;
                    16'hD5C0: data_out = 8'h95;
                    16'hD5C1: data_out = 8'h96;
                    16'hD5C2: data_out = 8'h97;
                    16'hD5C3: data_out = 8'h98;
                    16'hD5C4: data_out = 8'h99;
                    16'hD5C5: data_out = 8'h9A;
                    16'hD5C6: data_out = 8'h9B;
                    16'hD5C7: data_out = 8'h9C;
                    16'hD5C8: data_out = 8'h9D;
                    16'hD5C9: data_out = 8'h9E;
                    16'hD5CA: data_out = 8'h9F;
                    16'hD5CB: data_out = 8'hA0;
                    16'hD5CC: data_out = 8'hA1;
                    16'hD5CD: data_out = 8'hA2;
                    16'hD5CE: data_out = 8'hA3;
                    16'hD5CF: data_out = 8'hA4;
                    16'hD5D0: data_out = 8'hA5;
                    16'hD5D1: data_out = 8'hA6;
                    16'hD5D2: data_out = 8'hA7;
                    16'hD5D3: data_out = 8'hA8;
                    16'hD5D4: data_out = 8'hA9;
                    16'hD5D5: data_out = 8'hAA;
                    16'hD5D6: data_out = 8'hAB;
                    16'hD5D7: data_out = 8'hAC;
                    16'hD5D8: data_out = 8'hAD;
                    16'hD5D9: data_out = 8'hAE;
                    16'hD5DA: data_out = 8'hAF;
                    16'hD5DB: data_out = 8'hB0;
                    16'hD5DC: data_out = 8'hB1;
                    16'hD5DD: data_out = 8'hB2;
                    16'hD5DE: data_out = 8'hB3;
                    16'hD5DF: data_out = 8'hB4;
                    16'hD5E0: data_out = 8'hB5;
                    16'hD5E1: data_out = 8'hB6;
                    16'hD5E2: data_out = 8'hB7;
                    16'hD5E3: data_out = 8'hB8;
                    16'hD5E4: data_out = 8'hB9;
                    16'hD5E5: data_out = 8'hBA;
                    16'hD5E6: data_out = 8'hBB;
                    16'hD5E7: data_out = 8'hBC;
                    16'hD5E8: data_out = 8'hBD;
                    16'hD5E9: data_out = 8'hBE;
                    16'hD5EA: data_out = 8'hBF;
                    16'hD5EB: data_out = 8'hC0;
                    16'hD5EC: data_out = 8'hC1;
                    16'hD5ED: data_out = 8'hC2;
                    16'hD5EE: data_out = 8'hC3;
                    16'hD5EF: data_out = 8'hC4;
                    16'hD5F0: data_out = 8'hC5;
                    16'hD5F1: data_out = 8'hC6;
                    16'hD5F2: data_out = 8'hC7;
                    16'hD5F3: data_out = 8'hC8;
                    16'hD5F4: data_out = 8'hC9;
                    16'hD5F5: data_out = 8'hCA;
                    16'hD5F6: data_out = 8'hCB;
                    16'hD5F7: data_out = 8'hCC;
                    16'hD5F8: data_out = 8'hCD;
                    16'hD5F9: data_out = 8'hCE;
                    16'hD5FA: data_out = 8'hCF;
                    16'hD5FB: data_out = 8'hD0;
                    16'hD5FC: data_out = 8'hD1;
                    16'hD5FD: data_out = 8'hD2;
                    16'hD5FE: data_out = 8'hD3;
                    16'hD5FF: data_out = 8'hD4;
                    16'hD600: data_out = 8'hD6;
                    16'hD601: data_out = 8'hD5;
                    16'hD602: data_out = 8'hD4;
                    16'hD603: data_out = 8'hD3;
                    16'hD604: data_out = 8'hD2;
                    16'hD605: data_out = 8'hD1;
                    16'hD606: data_out = 8'hD0;
                    16'hD607: data_out = 8'hCF;
                    16'hD608: data_out = 8'hCE;
                    16'hD609: data_out = 8'hCD;
                    16'hD60A: data_out = 8'hCC;
                    16'hD60B: data_out = 8'hCB;
                    16'hD60C: data_out = 8'hCA;
                    16'hD60D: data_out = 8'hC9;
                    16'hD60E: data_out = 8'hC8;
                    16'hD60F: data_out = 8'hC7;
                    16'hD610: data_out = 8'hC6;
                    16'hD611: data_out = 8'hC5;
                    16'hD612: data_out = 8'hC4;
                    16'hD613: data_out = 8'hC3;
                    16'hD614: data_out = 8'hC2;
                    16'hD615: data_out = 8'hC1;
                    16'hD616: data_out = 8'hC0;
                    16'hD617: data_out = 8'hBF;
                    16'hD618: data_out = 8'hBE;
                    16'hD619: data_out = 8'hBD;
                    16'hD61A: data_out = 8'hBC;
                    16'hD61B: data_out = 8'hBB;
                    16'hD61C: data_out = 8'hBA;
                    16'hD61D: data_out = 8'hB9;
                    16'hD61E: data_out = 8'hB8;
                    16'hD61F: data_out = 8'hB7;
                    16'hD620: data_out = 8'hB6;
                    16'hD621: data_out = 8'hB5;
                    16'hD622: data_out = 8'hB4;
                    16'hD623: data_out = 8'hB3;
                    16'hD624: data_out = 8'hB2;
                    16'hD625: data_out = 8'hB1;
                    16'hD626: data_out = 8'hB0;
                    16'hD627: data_out = 8'hAF;
                    16'hD628: data_out = 8'hAE;
                    16'hD629: data_out = 8'hAD;
                    16'hD62A: data_out = 8'hAC;
                    16'hD62B: data_out = 8'hAB;
                    16'hD62C: data_out = 8'hAA;
                    16'hD62D: data_out = 8'hA9;
                    16'hD62E: data_out = 8'hA8;
                    16'hD62F: data_out = 8'hA7;
                    16'hD630: data_out = 8'hA6;
                    16'hD631: data_out = 8'hA5;
                    16'hD632: data_out = 8'hA4;
                    16'hD633: data_out = 8'hA3;
                    16'hD634: data_out = 8'hA2;
                    16'hD635: data_out = 8'hA1;
                    16'hD636: data_out = 8'hA0;
                    16'hD637: data_out = 8'h9F;
                    16'hD638: data_out = 8'h9E;
                    16'hD639: data_out = 8'h9D;
                    16'hD63A: data_out = 8'h9C;
                    16'hD63B: data_out = 8'h9B;
                    16'hD63C: data_out = 8'h9A;
                    16'hD63D: data_out = 8'h99;
                    16'hD63E: data_out = 8'h98;
                    16'hD63F: data_out = 8'h97;
                    16'hD640: data_out = 8'h96;
                    16'hD641: data_out = 8'h95;
                    16'hD642: data_out = 8'h94;
                    16'hD643: data_out = 8'h93;
                    16'hD644: data_out = 8'h92;
                    16'hD645: data_out = 8'h91;
                    16'hD646: data_out = 8'h90;
                    16'hD647: data_out = 8'h8F;
                    16'hD648: data_out = 8'h8E;
                    16'hD649: data_out = 8'h8D;
                    16'hD64A: data_out = 8'h8C;
                    16'hD64B: data_out = 8'h8B;
                    16'hD64C: data_out = 8'h8A;
                    16'hD64D: data_out = 8'h89;
                    16'hD64E: data_out = 8'h88;
                    16'hD64F: data_out = 8'h87;
                    16'hD650: data_out = 8'h86;
                    16'hD651: data_out = 8'h85;
                    16'hD652: data_out = 8'h84;
                    16'hD653: data_out = 8'h83;
                    16'hD654: data_out = 8'h82;
                    16'hD655: data_out = 8'h81;
                    16'hD656: data_out = 8'h0;
                    16'hD657: data_out = 8'h1;
                    16'hD658: data_out = 8'h2;
                    16'hD659: data_out = 8'h3;
                    16'hD65A: data_out = 8'h4;
                    16'hD65B: data_out = 8'h5;
                    16'hD65C: data_out = 8'h6;
                    16'hD65D: data_out = 8'h7;
                    16'hD65E: data_out = 8'h8;
                    16'hD65F: data_out = 8'h9;
                    16'hD660: data_out = 8'hA;
                    16'hD661: data_out = 8'hB;
                    16'hD662: data_out = 8'hC;
                    16'hD663: data_out = 8'hD;
                    16'hD664: data_out = 8'hE;
                    16'hD665: data_out = 8'hF;
                    16'hD666: data_out = 8'h10;
                    16'hD667: data_out = 8'h11;
                    16'hD668: data_out = 8'h12;
                    16'hD669: data_out = 8'h13;
                    16'hD66A: data_out = 8'h14;
                    16'hD66B: data_out = 8'h15;
                    16'hD66C: data_out = 8'h16;
                    16'hD66D: data_out = 8'h17;
                    16'hD66E: data_out = 8'h18;
                    16'hD66F: data_out = 8'h19;
                    16'hD670: data_out = 8'h1A;
                    16'hD671: data_out = 8'h1B;
                    16'hD672: data_out = 8'h1C;
                    16'hD673: data_out = 8'h1D;
                    16'hD674: data_out = 8'h1E;
                    16'hD675: data_out = 8'h1F;
                    16'hD676: data_out = 8'h20;
                    16'hD677: data_out = 8'h21;
                    16'hD678: data_out = 8'h22;
                    16'hD679: data_out = 8'h23;
                    16'hD67A: data_out = 8'h24;
                    16'hD67B: data_out = 8'h25;
                    16'hD67C: data_out = 8'h26;
                    16'hD67D: data_out = 8'h27;
                    16'hD67E: data_out = 8'h28;
                    16'hD67F: data_out = 8'h29;
                    16'hD680: data_out = 8'hD6;
                    16'hD681: data_out = 8'hD7;
                    16'hD682: data_out = 8'hD8;
                    16'hD683: data_out = 8'hD9;
                    16'hD684: data_out = 8'hDA;
                    16'hD685: data_out = 8'hDB;
                    16'hD686: data_out = 8'hDC;
                    16'hD687: data_out = 8'hDD;
                    16'hD688: data_out = 8'hDE;
                    16'hD689: data_out = 8'hDF;
                    16'hD68A: data_out = 8'hE0;
                    16'hD68B: data_out = 8'hE1;
                    16'hD68C: data_out = 8'hE2;
                    16'hD68D: data_out = 8'hE3;
                    16'hD68E: data_out = 8'hE4;
                    16'hD68F: data_out = 8'hE5;
                    16'hD690: data_out = 8'hE6;
                    16'hD691: data_out = 8'hE7;
                    16'hD692: data_out = 8'hE8;
                    16'hD693: data_out = 8'hE9;
                    16'hD694: data_out = 8'hEA;
                    16'hD695: data_out = 8'hEB;
                    16'hD696: data_out = 8'hEC;
                    16'hD697: data_out = 8'hED;
                    16'hD698: data_out = 8'hEE;
                    16'hD699: data_out = 8'hEF;
                    16'hD69A: data_out = 8'hF0;
                    16'hD69B: data_out = 8'hF1;
                    16'hD69C: data_out = 8'hF2;
                    16'hD69D: data_out = 8'hF3;
                    16'hD69E: data_out = 8'hF4;
                    16'hD69F: data_out = 8'hF5;
                    16'hD6A0: data_out = 8'hF6;
                    16'hD6A1: data_out = 8'hF7;
                    16'hD6A2: data_out = 8'hF8;
                    16'hD6A3: data_out = 8'hF9;
                    16'hD6A4: data_out = 8'hFA;
                    16'hD6A5: data_out = 8'hFB;
                    16'hD6A6: data_out = 8'hFC;
                    16'hD6A7: data_out = 8'hFD;
                    16'hD6A8: data_out = 8'hFE;
                    16'hD6A9: data_out = 8'hFF;
                    16'hD6AA: data_out = 8'h80;
                    16'hD6AB: data_out = 8'h81;
                    16'hD6AC: data_out = 8'h82;
                    16'hD6AD: data_out = 8'h83;
                    16'hD6AE: data_out = 8'h84;
                    16'hD6AF: data_out = 8'h85;
                    16'hD6B0: data_out = 8'h86;
                    16'hD6B1: data_out = 8'h87;
                    16'hD6B2: data_out = 8'h88;
                    16'hD6B3: data_out = 8'h89;
                    16'hD6B4: data_out = 8'h8A;
                    16'hD6B5: data_out = 8'h8B;
                    16'hD6B6: data_out = 8'h8C;
                    16'hD6B7: data_out = 8'h8D;
                    16'hD6B8: data_out = 8'h8E;
                    16'hD6B9: data_out = 8'h8F;
                    16'hD6BA: data_out = 8'h90;
                    16'hD6BB: data_out = 8'h91;
                    16'hD6BC: data_out = 8'h92;
                    16'hD6BD: data_out = 8'h93;
                    16'hD6BE: data_out = 8'h94;
                    16'hD6BF: data_out = 8'h95;
                    16'hD6C0: data_out = 8'h96;
                    16'hD6C1: data_out = 8'h97;
                    16'hD6C2: data_out = 8'h98;
                    16'hD6C3: data_out = 8'h99;
                    16'hD6C4: data_out = 8'h9A;
                    16'hD6C5: data_out = 8'h9B;
                    16'hD6C6: data_out = 8'h9C;
                    16'hD6C7: data_out = 8'h9D;
                    16'hD6C8: data_out = 8'h9E;
                    16'hD6C9: data_out = 8'h9F;
                    16'hD6CA: data_out = 8'hA0;
                    16'hD6CB: data_out = 8'hA1;
                    16'hD6CC: data_out = 8'hA2;
                    16'hD6CD: data_out = 8'hA3;
                    16'hD6CE: data_out = 8'hA4;
                    16'hD6CF: data_out = 8'hA5;
                    16'hD6D0: data_out = 8'hA6;
                    16'hD6D1: data_out = 8'hA7;
                    16'hD6D2: data_out = 8'hA8;
                    16'hD6D3: data_out = 8'hA9;
                    16'hD6D4: data_out = 8'hAA;
                    16'hD6D5: data_out = 8'hAB;
                    16'hD6D6: data_out = 8'hAC;
                    16'hD6D7: data_out = 8'hAD;
                    16'hD6D8: data_out = 8'hAE;
                    16'hD6D9: data_out = 8'hAF;
                    16'hD6DA: data_out = 8'hB0;
                    16'hD6DB: data_out = 8'hB1;
                    16'hD6DC: data_out = 8'hB2;
                    16'hD6DD: data_out = 8'hB3;
                    16'hD6DE: data_out = 8'hB4;
                    16'hD6DF: data_out = 8'hB5;
                    16'hD6E0: data_out = 8'hB6;
                    16'hD6E1: data_out = 8'hB7;
                    16'hD6E2: data_out = 8'hB8;
                    16'hD6E3: data_out = 8'hB9;
                    16'hD6E4: data_out = 8'hBA;
                    16'hD6E5: data_out = 8'hBB;
                    16'hD6E6: data_out = 8'hBC;
                    16'hD6E7: data_out = 8'hBD;
                    16'hD6E8: data_out = 8'hBE;
                    16'hD6E9: data_out = 8'hBF;
                    16'hD6EA: data_out = 8'hC0;
                    16'hD6EB: data_out = 8'hC1;
                    16'hD6EC: data_out = 8'hC2;
                    16'hD6ED: data_out = 8'hC3;
                    16'hD6EE: data_out = 8'hC4;
                    16'hD6EF: data_out = 8'hC5;
                    16'hD6F0: data_out = 8'hC6;
                    16'hD6F1: data_out = 8'hC7;
                    16'hD6F2: data_out = 8'hC8;
                    16'hD6F3: data_out = 8'hC9;
                    16'hD6F4: data_out = 8'hCA;
                    16'hD6F5: data_out = 8'hCB;
                    16'hD6F6: data_out = 8'hCC;
                    16'hD6F7: data_out = 8'hCD;
                    16'hD6F8: data_out = 8'hCE;
                    16'hD6F9: data_out = 8'hCF;
                    16'hD6FA: data_out = 8'hD0;
                    16'hD6FB: data_out = 8'hD1;
                    16'hD6FC: data_out = 8'hD2;
                    16'hD6FD: data_out = 8'hD3;
                    16'hD6FE: data_out = 8'hD4;
                    16'hD6FF: data_out = 8'hD5;
                    16'hD700: data_out = 8'hD7;
                    16'hD701: data_out = 8'hD6;
                    16'hD702: data_out = 8'hD5;
                    16'hD703: data_out = 8'hD4;
                    16'hD704: data_out = 8'hD3;
                    16'hD705: data_out = 8'hD2;
                    16'hD706: data_out = 8'hD1;
                    16'hD707: data_out = 8'hD0;
                    16'hD708: data_out = 8'hCF;
                    16'hD709: data_out = 8'hCE;
                    16'hD70A: data_out = 8'hCD;
                    16'hD70B: data_out = 8'hCC;
                    16'hD70C: data_out = 8'hCB;
                    16'hD70D: data_out = 8'hCA;
                    16'hD70E: data_out = 8'hC9;
                    16'hD70F: data_out = 8'hC8;
                    16'hD710: data_out = 8'hC7;
                    16'hD711: data_out = 8'hC6;
                    16'hD712: data_out = 8'hC5;
                    16'hD713: data_out = 8'hC4;
                    16'hD714: data_out = 8'hC3;
                    16'hD715: data_out = 8'hC2;
                    16'hD716: data_out = 8'hC1;
                    16'hD717: data_out = 8'hC0;
                    16'hD718: data_out = 8'hBF;
                    16'hD719: data_out = 8'hBE;
                    16'hD71A: data_out = 8'hBD;
                    16'hD71B: data_out = 8'hBC;
                    16'hD71C: data_out = 8'hBB;
                    16'hD71D: data_out = 8'hBA;
                    16'hD71E: data_out = 8'hB9;
                    16'hD71F: data_out = 8'hB8;
                    16'hD720: data_out = 8'hB7;
                    16'hD721: data_out = 8'hB6;
                    16'hD722: data_out = 8'hB5;
                    16'hD723: data_out = 8'hB4;
                    16'hD724: data_out = 8'hB3;
                    16'hD725: data_out = 8'hB2;
                    16'hD726: data_out = 8'hB1;
                    16'hD727: data_out = 8'hB0;
                    16'hD728: data_out = 8'hAF;
                    16'hD729: data_out = 8'hAE;
                    16'hD72A: data_out = 8'hAD;
                    16'hD72B: data_out = 8'hAC;
                    16'hD72C: data_out = 8'hAB;
                    16'hD72D: data_out = 8'hAA;
                    16'hD72E: data_out = 8'hA9;
                    16'hD72F: data_out = 8'hA8;
                    16'hD730: data_out = 8'hA7;
                    16'hD731: data_out = 8'hA6;
                    16'hD732: data_out = 8'hA5;
                    16'hD733: data_out = 8'hA4;
                    16'hD734: data_out = 8'hA3;
                    16'hD735: data_out = 8'hA2;
                    16'hD736: data_out = 8'hA1;
                    16'hD737: data_out = 8'hA0;
                    16'hD738: data_out = 8'h9F;
                    16'hD739: data_out = 8'h9E;
                    16'hD73A: data_out = 8'h9D;
                    16'hD73B: data_out = 8'h9C;
                    16'hD73C: data_out = 8'h9B;
                    16'hD73D: data_out = 8'h9A;
                    16'hD73E: data_out = 8'h99;
                    16'hD73F: data_out = 8'h98;
                    16'hD740: data_out = 8'h97;
                    16'hD741: data_out = 8'h96;
                    16'hD742: data_out = 8'h95;
                    16'hD743: data_out = 8'h94;
                    16'hD744: data_out = 8'h93;
                    16'hD745: data_out = 8'h92;
                    16'hD746: data_out = 8'h91;
                    16'hD747: data_out = 8'h90;
                    16'hD748: data_out = 8'h8F;
                    16'hD749: data_out = 8'h8E;
                    16'hD74A: data_out = 8'h8D;
                    16'hD74B: data_out = 8'h8C;
                    16'hD74C: data_out = 8'h8B;
                    16'hD74D: data_out = 8'h8A;
                    16'hD74E: data_out = 8'h89;
                    16'hD74F: data_out = 8'h88;
                    16'hD750: data_out = 8'h87;
                    16'hD751: data_out = 8'h86;
                    16'hD752: data_out = 8'h85;
                    16'hD753: data_out = 8'h84;
                    16'hD754: data_out = 8'h83;
                    16'hD755: data_out = 8'h82;
                    16'hD756: data_out = 8'h81;
                    16'hD757: data_out = 8'h0;
                    16'hD758: data_out = 8'h1;
                    16'hD759: data_out = 8'h2;
                    16'hD75A: data_out = 8'h3;
                    16'hD75B: data_out = 8'h4;
                    16'hD75C: data_out = 8'h5;
                    16'hD75D: data_out = 8'h6;
                    16'hD75E: data_out = 8'h7;
                    16'hD75F: data_out = 8'h8;
                    16'hD760: data_out = 8'h9;
                    16'hD761: data_out = 8'hA;
                    16'hD762: data_out = 8'hB;
                    16'hD763: data_out = 8'hC;
                    16'hD764: data_out = 8'hD;
                    16'hD765: data_out = 8'hE;
                    16'hD766: data_out = 8'hF;
                    16'hD767: data_out = 8'h10;
                    16'hD768: data_out = 8'h11;
                    16'hD769: data_out = 8'h12;
                    16'hD76A: data_out = 8'h13;
                    16'hD76B: data_out = 8'h14;
                    16'hD76C: data_out = 8'h15;
                    16'hD76D: data_out = 8'h16;
                    16'hD76E: data_out = 8'h17;
                    16'hD76F: data_out = 8'h18;
                    16'hD770: data_out = 8'h19;
                    16'hD771: data_out = 8'h1A;
                    16'hD772: data_out = 8'h1B;
                    16'hD773: data_out = 8'h1C;
                    16'hD774: data_out = 8'h1D;
                    16'hD775: data_out = 8'h1E;
                    16'hD776: data_out = 8'h1F;
                    16'hD777: data_out = 8'h20;
                    16'hD778: data_out = 8'h21;
                    16'hD779: data_out = 8'h22;
                    16'hD77A: data_out = 8'h23;
                    16'hD77B: data_out = 8'h24;
                    16'hD77C: data_out = 8'h25;
                    16'hD77D: data_out = 8'h26;
                    16'hD77E: data_out = 8'h27;
                    16'hD77F: data_out = 8'h28;
                    16'hD780: data_out = 8'hD7;
                    16'hD781: data_out = 8'hD8;
                    16'hD782: data_out = 8'hD9;
                    16'hD783: data_out = 8'hDA;
                    16'hD784: data_out = 8'hDB;
                    16'hD785: data_out = 8'hDC;
                    16'hD786: data_out = 8'hDD;
                    16'hD787: data_out = 8'hDE;
                    16'hD788: data_out = 8'hDF;
                    16'hD789: data_out = 8'hE0;
                    16'hD78A: data_out = 8'hE1;
                    16'hD78B: data_out = 8'hE2;
                    16'hD78C: data_out = 8'hE3;
                    16'hD78D: data_out = 8'hE4;
                    16'hD78E: data_out = 8'hE5;
                    16'hD78F: data_out = 8'hE6;
                    16'hD790: data_out = 8'hE7;
                    16'hD791: data_out = 8'hE8;
                    16'hD792: data_out = 8'hE9;
                    16'hD793: data_out = 8'hEA;
                    16'hD794: data_out = 8'hEB;
                    16'hD795: data_out = 8'hEC;
                    16'hD796: data_out = 8'hED;
                    16'hD797: data_out = 8'hEE;
                    16'hD798: data_out = 8'hEF;
                    16'hD799: data_out = 8'hF0;
                    16'hD79A: data_out = 8'hF1;
                    16'hD79B: data_out = 8'hF2;
                    16'hD79C: data_out = 8'hF3;
                    16'hD79D: data_out = 8'hF4;
                    16'hD79E: data_out = 8'hF5;
                    16'hD79F: data_out = 8'hF6;
                    16'hD7A0: data_out = 8'hF7;
                    16'hD7A1: data_out = 8'hF8;
                    16'hD7A2: data_out = 8'hF9;
                    16'hD7A3: data_out = 8'hFA;
                    16'hD7A4: data_out = 8'hFB;
                    16'hD7A5: data_out = 8'hFC;
                    16'hD7A6: data_out = 8'hFD;
                    16'hD7A7: data_out = 8'hFE;
                    16'hD7A8: data_out = 8'hFF;
                    16'hD7A9: data_out = 8'h80;
                    16'hD7AA: data_out = 8'h81;
                    16'hD7AB: data_out = 8'h82;
                    16'hD7AC: data_out = 8'h83;
                    16'hD7AD: data_out = 8'h84;
                    16'hD7AE: data_out = 8'h85;
                    16'hD7AF: data_out = 8'h86;
                    16'hD7B0: data_out = 8'h87;
                    16'hD7B1: data_out = 8'h88;
                    16'hD7B2: data_out = 8'h89;
                    16'hD7B3: data_out = 8'h8A;
                    16'hD7B4: data_out = 8'h8B;
                    16'hD7B5: data_out = 8'h8C;
                    16'hD7B6: data_out = 8'h8D;
                    16'hD7B7: data_out = 8'h8E;
                    16'hD7B8: data_out = 8'h8F;
                    16'hD7B9: data_out = 8'h90;
                    16'hD7BA: data_out = 8'h91;
                    16'hD7BB: data_out = 8'h92;
                    16'hD7BC: data_out = 8'h93;
                    16'hD7BD: data_out = 8'h94;
                    16'hD7BE: data_out = 8'h95;
                    16'hD7BF: data_out = 8'h96;
                    16'hD7C0: data_out = 8'h97;
                    16'hD7C1: data_out = 8'h98;
                    16'hD7C2: data_out = 8'h99;
                    16'hD7C3: data_out = 8'h9A;
                    16'hD7C4: data_out = 8'h9B;
                    16'hD7C5: data_out = 8'h9C;
                    16'hD7C6: data_out = 8'h9D;
                    16'hD7C7: data_out = 8'h9E;
                    16'hD7C8: data_out = 8'h9F;
                    16'hD7C9: data_out = 8'hA0;
                    16'hD7CA: data_out = 8'hA1;
                    16'hD7CB: data_out = 8'hA2;
                    16'hD7CC: data_out = 8'hA3;
                    16'hD7CD: data_out = 8'hA4;
                    16'hD7CE: data_out = 8'hA5;
                    16'hD7CF: data_out = 8'hA6;
                    16'hD7D0: data_out = 8'hA7;
                    16'hD7D1: data_out = 8'hA8;
                    16'hD7D2: data_out = 8'hA9;
                    16'hD7D3: data_out = 8'hAA;
                    16'hD7D4: data_out = 8'hAB;
                    16'hD7D5: data_out = 8'hAC;
                    16'hD7D6: data_out = 8'hAD;
                    16'hD7D7: data_out = 8'hAE;
                    16'hD7D8: data_out = 8'hAF;
                    16'hD7D9: data_out = 8'hB0;
                    16'hD7DA: data_out = 8'hB1;
                    16'hD7DB: data_out = 8'hB2;
                    16'hD7DC: data_out = 8'hB3;
                    16'hD7DD: data_out = 8'hB4;
                    16'hD7DE: data_out = 8'hB5;
                    16'hD7DF: data_out = 8'hB6;
                    16'hD7E0: data_out = 8'hB7;
                    16'hD7E1: data_out = 8'hB8;
                    16'hD7E2: data_out = 8'hB9;
                    16'hD7E3: data_out = 8'hBA;
                    16'hD7E4: data_out = 8'hBB;
                    16'hD7E5: data_out = 8'hBC;
                    16'hD7E6: data_out = 8'hBD;
                    16'hD7E7: data_out = 8'hBE;
                    16'hD7E8: data_out = 8'hBF;
                    16'hD7E9: data_out = 8'hC0;
                    16'hD7EA: data_out = 8'hC1;
                    16'hD7EB: data_out = 8'hC2;
                    16'hD7EC: data_out = 8'hC3;
                    16'hD7ED: data_out = 8'hC4;
                    16'hD7EE: data_out = 8'hC5;
                    16'hD7EF: data_out = 8'hC6;
                    16'hD7F0: data_out = 8'hC7;
                    16'hD7F1: data_out = 8'hC8;
                    16'hD7F2: data_out = 8'hC9;
                    16'hD7F3: data_out = 8'hCA;
                    16'hD7F4: data_out = 8'hCB;
                    16'hD7F5: data_out = 8'hCC;
                    16'hD7F6: data_out = 8'hCD;
                    16'hD7F7: data_out = 8'hCE;
                    16'hD7F8: data_out = 8'hCF;
                    16'hD7F9: data_out = 8'hD0;
                    16'hD7FA: data_out = 8'hD1;
                    16'hD7FB: data_out = 8'hD2;
                    16'hD7FC: data_out = 8'hD3;
                    16'hD7FD: data_out = 8'hD4;
                    16'hD7FE: data_out = 8'hD5;
                    16'hD7FF: data_out = 8'hD6;
                    16'hD800: data_out = 8'hD8;
                    16'hD801: data_out = 8'hD7;
                    16'hD802: data_out = 8'hD6;
                    16'hD803: data_out = 8'hD5;
                    16'hD804: data_out = 8'hD4;
                    16'hD805: data_out = 8'hD3;
                    16'hD806: data_out = 8'hD2;
                    16'hD807: data_out = 8'hD1;
                    16'hD808: data_out = 8'hD0;
                    16'hD809: data_out = 8'hCF;
                    16'hD80A: data_out = 8'hCE;
                    16'hD80B: data_out = 8'hCD;
                    16'hD80C: data_out = 8'hCC;
                    16'hD80D: data_out = 8'hCB;
                    16'hD80E: data_out = 8'hCA;
                    16'hD80F: data_out = 8'hC9;
                    16'hD810: data_out = 8'hC8;
                    16'hD811: data_out = 8'hC7;
                    16'hD812: data_out = 8'hC6;
                    16'hD813: data_out = 8'hC5;
                    16'hD814: data_out = 8'hC4;
                    16'hD815: data_out = 8'hC3;
                    16'hD816: data_out = 8'hC2;
                    16'hD817: data_out = 8'hC1;
                    16'hD818: data_out = 8'hC0;
                    16'hD819: data_out = 8'hBF;
                    16'hD81A: data_out = 8'hBE;
                    16'hD81B: data_out = 8'hBD;
                    16'hD81C: data_out = 8'hBC;
                    16'hD81D: data_out = 8'hBB;
                    16'hD81E: data_out = 8'hBA;
                    16'hD81F: data_out = 8'hB9;
                    16'hD820: data_out = 8'hB8;
                    16'hD821: data_out = 8'hB7;
                    16'hD822: data_out = 8'hB6;
                    16'hD823: data_out = 8'hB5;
                    16'hD824: data_out = 8'hB4;
                    16'hD825: data_out = 8'hB3;
                    16'hD826: data_out = 8'hB2;
                    16'hD827: data_out = 8'hB1;
                    16'hD828: data_out = 8'hB0;
                    16'hD829: data_out = 8'hAF;
                    16'hD82A: data_out = 8'hAE;
                    16'hD82B: data_out = 8'hAD;
                    16'hD82C: data_out = 8'hAC;
                    16'hD82D: data_out = 8'hAB;
                    16'hD82E: data_out = 8'hAA;
                    16'hD82F: data_out = 8'hA9;
                    16'hD830: data_out = 8'hA8;
                    16'hD831: data_out = 8'hA7;
                    16'hD832: data_out = 8'hA6;
                    16'hD833: data_out = 8'hA5;
                    16'hD834: data_out = 8'hA4;
                    16'hD835: data_out = 8'hA3;
                    16'hD836: data_out = 8'hA2;
                    16'hD837: data_out = 8'hA1;
                    16'hD838: data_out = 8'hA0;
                    16'hD839: data_out = 8'h9F;
                    16'hD83A: data_out = 8'h9E;
                    16'hD83B: data_out = 8'h9D;
                    16'hD83C: data_out = 8'h9C;
                    16'hD83D: data_out = 8'h9B;
                    16'hD83E: data_out = 8'h9A;
                    16'hD83F: data_out = 8'h99;
                    16'hD840: data_out = 8'h98;
                    16'hD841: data_out = 8'h97;
                    16'hD842: data_out = 8'h96;
                    16'hD843: data_out = 8'h95;
                    16'hD844: data_out = 8'h94;
                    16'hD845: data_out = 8'h93;
                    16'hD846: data_out = 8'h92;
                    16'hD847: data_out = 8'h91;
                    16'hD848: data_out = 8'h90;
                    16'hD849: data_out = 8'h8F;
                    16'hD84A: data_out = 8'h8E;
                    16'hD84B: data_out = 8'h8D;
                    16'hD84C: data_out = 8'h8C;
                    16'hD84D: data_out = 8'h8B;
                    16'hD84E: data_out = 8'h8A;
                    16'hD84F: data_out = 8'h89;
                    16'hD850: data_out = 8'h88;
                    16'hD851: data_out = 8'h87;
                    16'hD852: data_out = 8'h86;
                    16'hD853: data_out = 8'h85;
                    16'hD854: data_out = 8'h84;
                    16'hD855: data_out = 8'h83;
                    16'hD856: data_out = 8'h82;
                    16'hD857: data_out = 8'h81;
                    16'hD858: data_out = 8'h0;
                    16'hD859: data_out = 8'h1;
                    16'hD85A: data_out = 8'h2;
                    16'hD85B: data_out = 8'h3;
                    16'hD85C: data_out = 8'h4;
                    16'hD85D: data_out = 8'h5;
                    16'hD85E: data_out = 8'h6;
                    16'hD85F: data_out = 8'h7;
                    16'hD860: data_out = 8'h8;
                    16'hD861: data_out = 8'h9;
                    16'hD862: data_out = 8'hA;
                    16'hD863: data_out = 8'hB;
                    16'hD864: data_out = 8'hC;
                    16'hD865: data_out = 8'hD;
                    16'hD866: data_out = 8'hE;
                    16'hD867: data_out = 8'hF;
                    16'hD868: data_out = 8'h10;
                    16'hD869: data_out = 8'h11;
                    16'hD86A: data_out = 8'h12;
                    16'hD86B: data_out = 8'h13;
                    16'hD86C: data_out = 8'h14;
                    16'hD86D: data_out = 8'h15;
                    16'hD86E: data_out = 8'h16;
                    16'hD86F: data_out = 8'h17;
                    16'hD870: data_out = 8'h18;
                    16'hD871: data_out = 8'h19;
                    16'hD872: data_out = 8'h1A;
                    16'hD873: data_out = 8'h1B;
                    16'hD874: data_out = 8'h1C;
                    16'hD875: data_out = 8'h1D;
                    16'hD876: data_out = 8'h1E;
                    16'hD877: data_out = 8'h1F;
                    16'hD878: data_out = 8'h20;
                    16'hD879: data_out = 8'h21;
                    16'hD87A: data_out = 8'h22;
                    16'hD87B: data_out = 8'h23;
                    16'hD87C: data_out = 8'h24;
                    16'hD87D: data_out = 8'h25;
                    16'hD87E: data_out = 8'h26;
                    16'hD87F: data_out = 8'h27;
                    16'hD880: data_out = 8'hD8;
                    16'hD881: data_out = 8'hD9;
                    16'hD882: data_out = 8'hDA;
                    16'hD883: data_out = 8'hDB;
                    16'hD884: data_out = 8'hDC;
                    16'hD885: data_out = 8'hDD;
                    16'hD886: data_out = 8'hDE;
                    16'hD887: data_out = 8'hDF;
                    16'hD888: data_out = 8'hE0;
                    16'hD889: data_out = 8'hE1;
                    16'hD88A: data_out = 8'hE2;
                    16'hD88B: data_out = 8'hE3;
                    16'hD88C: data_out = 8'hE4;
                    16'hD88D: data_out = 8'hE5;
                    16'hD88E: data_out = 8'hE6;
                    16'hD88F: data_out = 8'hE7;
                    16'hD890: data_out = 8'hE8;
                    16'hD891: data_out = 8'hE9;
                    16'hD892: data_out = 8'hEA;
                    16'hD893: data_out = 8'hEB;
                    16'hD894: data_out = 8'hEC;
                    16'hD895: data_out = 8'hED;
                    16'hD896: data_out = 8'hEE;
                    16'hD897: data_out = 8'hEF;
                    16'hD898: data_out = 8'hF0;
                    16'hD899: data_out = 8'hF1;
                    16'hD89A: data_out = 8'hF2;
                    16'hD89B: data_out = 8'hF3;
                    16'hD89C: data_out = 8'hF4;
                    16'hD89D: data_out = 8'hF5;
                    16'hD89E: data_out = 8'hF6;
                    16'hD89F: data_out = 8'hF7;
                    16'hD8A0: data_out = 8'hF8;
                    16'hD8A1: data_out = 8'hF9;
                    16'hD8A2: data_out = 8'hFA;
                    16'hD8A3: data_out = 8'hFB;
                    16'hD8A4: data_out = 8'hFC;
                    16'hD8A5: data_out = 8'hFD;
                    16'hD8A6: data_out = 8'hFE;
                    16'hD8A7: data_out = 8'hFF;
                    16'hD8A8: data_out = 8'h80;
                    16'hD8A9: data_out = 8'h81;
                    16'hD8AA: data_out = 8'h82;
                    16'hD8AB: data_out = 8'h83;
                    16'hD8AC: data_out = 8'h84;
                    16'hD8AD: data_out = 8'h85;
                    16'hD8AE: data_out = 8'h86;
                    16'hD8AF: data_out = 8'h87;
                    16'hD8B0: data_out = 8'h88;
                    16'hD8B1: data_out = 8'h89;
                    16'hD8B2: data_out = 8'h8A;
                    16'hD8B3: data_out = 8'h8B;
                    16'hD8B4: data_out = 8'h8C;
                    16'hD8B5: data_out = 8'h8D;
                    16'hD8B6: data_out = 8'h8E;
                    16'hD8B7: data_out = 8'h8F;
                    16'hD8B8: data_out = 8'h90;
                    16'hD8B9: data_out = 8'h91;
                    16'hD8BA: data_out = 8'h92;
                    16'hD8BB: data_out = 8'h93;
                    16'hD8BC: data_out = 8'h94;
                    16'hD8BD: data_out = 8'h95;
                    16'hD8BE: data_out = 8'h96;
                    16'hD8BF: data_out = 8'h97;
                    16'hD8C0: data_out = 8'h98;
                    16'hD8C1: data_out = 8'h99;
                    16'hD8C2: data_out = 8'h9A;
                    16'hD8C3: data_out = 8'h9B;
                    16'hD8C4: data_out = 8'h9C;
                    16'hD8C5: data_out = 8'h9D;
                    16'hD8C6: data_out = 8'h9E;
                    16'hD8C7: data_out = 8'h9F;
                    16'hD8C8: data_out = 8'hA0;
                    16'hD8C9: data_out = 8'hA1;
                    16'hD8CA: data_out = 8'hA2;
                    16'hD8CB: data_out = 8'hA3;
                    16'hD8CC: data_out = 8'hA4;
                    16'hD8CD: data_out = 8'hA5;
                    16'hD8CE: data_out = 8'hA6;
                    16'hD8CF: data_out = 8'hA7;
                    16'hD8D0: data_out = 8'hA8;
                    16'hD8D1: data_out = 8'hA9;
                    16'hD8D2: data_out = 8'hAA;
                    16'hD8D3: data_out = 8'hAB;
                    16'hD8D4: data_out = 8'hAC;
                    16'hD8D5: data_out = 8'hAD;
                    16'hD8D6: data_out = 8'hAE;
                    16'hD8D7: data_out = 8'hAF;
                    16'hD8D8: data_out = 8'hB0;
                    16'hD8D9: data_out = 8'hB1;
                    16'hD8DA: data_out = 8'hB2;
                    16'hD8DB: data_out = 8'hB3;
                    16'hD8DC: data_out = 8'hB4;
                    16'hD8DD: data_out = 8'hB5;
                    16'hD8DE: data_out = 8'hB6;
                    16'hD8DF: data_out = 8'hB7;
                    16'hD8E0: data_out = 8'hB8;
                    16'hD8E1: data_out = 8'hB9;
                    16'hD8E2: data_out = 8'hBA;
                    16'hD8E3: data_out = 8'hBB;
                    16'hD8E4: data_out = 8'hBC;
                    16'hD8E5: data_out = 8'hBD;
                    16'hD8E6: data_out = 8'hBE;
                    16'hD8E7: data_out = 8'hBF;
                    16'hD8E8: data_out = 8'hC0;
                    16'hD8E9: data_out = 8'hC1;
                    16'hD8EA: data_out = 8'hC2;
                    16'hD8EB: data_out = 8'hC3;
                    16'hD8EC: data_out = 8'hC4;
                    16'hD8ED: data_out = 8'hC5;
                    16'hD8EE: data_out = 8'hC6;
                    16'hD8EF: data_out = 8'hC7;
                    16'hD8F0: data_out = 8'hC8;
                    16'hD8F1: data_out = 8'hC9;
                    16'hD8F2: data_out = 8'hCA;
                    16'hD8F3: data_out = 8'hCB;
                    16'hD8F4: data_out = 8'hCC;
                    16'hD8F5: data_out = 8'hCD;
                    16'hD8F6: data_out = 8'hCE;
                    16'hD8F7: data_out = 8'hCF;
                    16'hD8F8: data_out = 8'hD0;
                    16'hD8F9: data_out = 8'hD1;
                    16'hD8FA: data_out = 8'hD2;
                    16'hD8FB: data_out = 8'hD3;
                    16'hD8FC: data_out = 8'hD4;
                    16'hD8FD: data_out = 8'hD5;
                    16'hD8FE: data_out = 8'hD6;
                    16'hD8FF: data_out = 8'hD7;
                    16'hD900: data_out = 8'hD9;
                    16'hD901: data_out = 8'hD8;
                    16'hD902: data_out = 8'hD7;
                    16'hD903: data_out = 8'hD6;
                    16'hD904: data_out = 8'hD5;
                    16'hD905: data_out = 8'hD4;
                    16'hD906: data_out = 8'hD3;
                    16'hD907: data_out = 8'hD2;
                    16'hD908: data_out = 8'hD1;
                    16'hD909: data_out = 8'hD0;
                    16'hD90A: data_out = 8'hCF;
                    16'hD90B: data_out = 8'hCE;
                    16'hD90C: data_out = 8'hCD;
                    16'hD90D: data_out = 8'hCC;
                    16'hD90E: data_out = 8'hCB;
                    16'hD90F: data_out = 8'hCA;
                    16'hD910: data_out = 8'hC9;
                    16'hD911: data_out = 8'hC8;
                    16'hD912: data_out = 8'hC7;
                    16'hD913: data_out = 8'hC6;
                    16'hD914: data_out = 8'hC5;
                    16'hD915: data_out = 8'hC4;
                    16'hD916: data_out = 8'hC3;
                    16'hD917: data_out = 8'hC2;
                    16'hD918: data_out = 8'hC1;
                    16'hD919: data_out = 8'hC0;
                    16'hD91A: data_out = 8'hBF;
                    16'hD91B: data_out = 8'hBE;
                    16'hD91C: data_out = 8'hBD;
                    16'hD91D: data_out = 8'hBC;
                    16'hD91E: data_out = 8'hBB;
                    16'hD91F: data_out = 8'hBA;
                    16'hD920: data_out = 8'hB9;
                    16'hD921: data_out = 8'hB8;
                    16'hD922: data_out = 8'hB7;
                    16'hD923: data_out = 8'hB6;
                    16'hD924: data_out = 8'hB5;
                    16'hD925: data_out = 8'hB4;
                    16'hD926: data_out = 8'hB3;
                    16'hD927: data_out = 8'hB2;
                    16'hD928: data_out = 8'hB1;
                    16'hD929: data_out = 8'hB0;
                    16'hD92A: data_out = 8'hAF;
                    16'hD92B: data_out = 8'hAE;
                    16'hD92C: data_out = 8'hAD;
                    16'hD92D: data_out = 8'hAC;
                    16'hD92E: data_out = 8'hAB;
                    16'hD92F: data_out = 8'hAA;
                    16'hD930: data_out = 8'hA9;
                    16'hD931: data_out = 8'hA8;
                    16'hD932: data_out = 8'hA7;
                    16'hD933: data_out = 8'hA6;
                    16'hD934: data_out = 8'hA5;
                    16'hD935: data_out = 8'hA4;
                    16'hD936: data_out = 8'hA3;
                    16'hD937: data_out = 8'hA2;
                    16'hD938: data_out = 8'hA1;
                    16'hD939: data_out = 8'hA0;
                    16'hD93A: data_out = 8'h9F;
                    16'hD93B: data_out = 8'h9E;
                    16'hD93C: data_out = 8'h9D;
                    16'hD93D: data_out = 8'h9C;
                    16'hD93E: data_out = 8'h9B;
                    16'hD93F: data_out = 8'h9A;
                    16'hD940: data_out = 8'h99;
                    16'hD941: data_out = 8'h98;
                    16'hD942: data_out = 8'h97;
                    16'hD943: data_out = 8'h96;
                    16'hD944: data_out = 8'h95;
                    16'hD945: data_out = 8'h94;
                    16'hD946: data_out = 8'h93;
                    16'hD947: data_out = 8'h92;
                    16'hD948: data_out = 8'h91;
                    16'hD949: data_out = 8'h90;
                    16'hD94A: data_out = 8'h8F;
                    16'hD94B: data_out = 8'h8E;
                    16'hD94C: data_out = 8'h8D;
                    16'hD94D: data_out = 8'h8C;
                    16'hD94E: data_out = 8'h8B;
                    16'hD94F: data_out = 8'h8A;
                    16'hD950: data_out = 8'h89;
                    16'hD951: data_out = 8'h88;
                    16'hD952: data_out = 8'h87;
                    16'hD953: data_out = 8'h86;
                    16'hD954: data_out = 8'h85;
                    16'hD955: data_out = 8'h84;
                    16'hD956: data_out = 8'h83;
                    16'hD957: data_out = 8'h82;
                    16'hD958: data_out = 8'h81;
                    16'hD959: data_out = 8'h0;
                    16'hD95A: data_out = 8'h1;
                    16'hD95B: data_out = 8'h2;
                    16'hD95C: data_out = 8'h3;
                    16'hD95D: data_out = 8'h4;
                    16'hD95E: data_out = 8'h5;
                    16'hD95F: data_out = 8'h6;
                    16'hD960: data_out = 8'h7;
                    16'hD961: data_out = 8'h8;
                    16'hD962: data_out = 8'h9;
                    16'hD963: data_out = 8'hA;
                    16'hD964: data_out = 8'hB;
                    16'hD965: data_out = 8'hC;
                    16'hD966: data_out = 8'hD;
                    16'hD967: data_out = 8'hE;
                    16'hD968: data_out = 8'hF;
                    16'hD969: data_out = 8'h10;
                    16'hD96A: data_out = 8'h11;
                    16'hD96B: data_out = 8'h12;
                    16'hD96C: data_out = 8'h13;
                    16'hD96D: data_out = 8'h14;
                    16'hD96E: data_out = 8'h15;
                    16'hD96F: data_out = 8'h16;
                    16'hD970: data_out = 8'h17;
                    16'hD971: data_out = 8'h18;
                    16'hD972: data_out = 8'h19;
                    16'hD973: data_out = 8'h1A;
                    16'hD974: data_out = 8'h1B;
                    16'hD975: data_out = 8'h1C;
                    16'hD976: data_out = 8'h1D;
                    16'hD977: data_out = 8'h1E;
                    16'hD978: data_out = 8'h1F;
                    16'hD979: data_out = 8'h20;
                    16'hD97A: data_out = 8'h21;
                    16'hD97B: data_out = 8'h22;
                    16'hD97C: data_out = 8'h23;
                    16'hD97D: data_out = 8'h24;
                    16'hD97E: data_out = 8'h25;
                    16'hD97F: data_out = 8'h26;
                    16'hD980: data_out = 8'hD9;
                    16'hD981: data_out = 8'hDA;
                    16'hD982: data_out = 8'hDB;
                    16'hD983: data_out = 8'hDC;
                    16'hD984: data_out = 8'hDD;
                    16'hD985: data_out = 8'hDE;
                    16'hD986: data_out = 8'hDF;
                    16'hD987: data_out = 8'hE0;
                    16'hD988: data_out = 8'hE1;
                    16'hD989: data_out = 8'hE2;
                    16'hD98A: data_out = 8'hE3;
                    16'hD98B: data_out = 8'hE4;
                    16'hD98C: data_out = 8'hE5;
                    16'hD98D: data_out = 8'hE6;
                    16'hD98E: data_out = 8'hE7;
                    16'hD98F: data_out = 8'hE8;
                    16'hD990: data_out = 8'hE9;
                    16'hD991: data_out = 8'hEA;
                    16'hD992: data_out = 8'hEB;
                    16'hD993: data_out = 8'hEC;
                    16'hD994: data_out = 8'hED;
                    16'hD995: data_out = 8'hEE;
                    16'hD996: data_out = 8'hEF;
                    16'hD997: data_out = 8'hF0;
                    16'hD998: data_out = 8'hF1;
                    16'hD999: data_out = 8'hF2;
                    16'hD99A: data_out = 8'hF3;
                    16'hD99B: data_out = 8'hF4;
                    16'hD99C: data_out = 8'hF5;
                    16'hD99D: data_out = 8'hF6;
                    16'hD99E: data_out = 8'hF7;
                    16'hD99F: data_out = 8'hF8;
                    16'hD9A0: data_out = 8'hF9;
                    16'hD9A1: data_out = 8'hFA;
                    16'hD9A2: data_out = 8'hFB;
                    16'hD9A3: data_out = 8'hFC;
                    16'hD9A4: data_out = 8'hFD;
                    16'hD9A5: data_out = 8'hFE;
                    16'hD9A6: data_out = 8'hFF;
                    16'hD9A7: data_out = 8'h80;
                    16'hD9A8: data_out = 8'h81;
                    16'hD9A9: data_out = 8'h82;
                    16'hD9AA: data_out = 8'h83;
                    16'hD9AB: data_out = 8'h84;
                    16'hD9AC: data_out = 8'h85;
                    16'hD9AD: data_out = 8'h86;
                    16'hD9AE: data_out = 8'h87;
                    16'hD9AF: data_out = 8'h88;
                    16'hD9B0: data_out = 8'h89;
                    16'hD9B1: data_out = 8'h8A;
                    16'hD9B2: data_out = 8'h8B;
                    16'hD9B3: data_out = 8'h8C;
                    16'hD9B4: data_out = 8'h8D;
                    16'hD9B5: data_out = 8'h8E;
                    16'hD9B6: data_out = 8'h8F;
                    16'hD9B7: data_out = 8'h90;
                    16'hD9B8: data_out = 8'h91;
                    16'hD9B9: data_out = 8'h92;
                    16'hD9BA: data_out = 8'h93;
                    16'hD9BB: data_out = 8'h94;
                    16'hD9BC: data_out = 8'h95;
                    16'hD9BD: data_out = 8'h96;
                    16'hD9BE: data_out = 8'h97;
                    16'hD9BF: data_out = 8'h98;
                    16'hD9C0: data_out = 8'h99;
                    16'hD9C1: data_out = 8'h9A;
                    16'hD9C2: data_out = 8'h9B;
                    16'hD9C3: data_out = 8'h9C;
                    16'hD9C4: data_out = 8'h9D;
                    16'hD9C5: data_out = 8'h9E;
                    16'hD9C6: data_out = 8'h9F;
                    16'hD9C7: data_out = 8'hA0;
                    16'hD9C8: data_out = 8'hA1;
                    16'hD9C9: data_out = 8'hA2;
                    16'hD9CA: data_out = 8'hA3;
                    16'hD9CB: data_out = 8'hA4;
                    16'hD9CC: data_out = 8'hA5;
                    16'hD9CD: data_out = 8'hA6;
                    16'hD9CE: data_out = 8'hA7;
                    16'hD9CF: data_out = 8'hA8;
                    16'hD9D0: data_out = 8'hA9;
                    16'hD9D1: data_out = 8'hAA;
                    16'hD9D2: data_out = 8'hAB;
                    16'hD9D3: data_out = 8'hAC;
                    16'hD9D4: data_out = 8'hAD;
                    16'hD9D5: data_out = 8'hAE;
                    16'hD9D6: data_out = 8'hAF;
                    16'hD9D7: data_out = 8'hB0;
                    16'hD9D8: data_out = 8'hB1;
                    16'hD9D9: data_out = 8'hB2;
                    16'hD9DA: data_out = 8'hB3;
                    16'hD9DB: data_out = 8'hB4;
                    16'hD9DC: data_out = 8'hB5;
                    16'hD9DD: data_out = 8'hB6;
                    16'hD9DE: data_out = 8'hB7;
                    16'hD9DF: data_out = 8'hB8;
                    16'hD9E0: data_out = 8'hB9;
                    16'hD9E1: data_out = 8'hBA;
                    16'hD9E2: data_out = 8'hBB;
                    16'hD9E3: data_out = 8'hBC;
                    16'hD9E4: data_out = 8'hBD;
                    16'hD9E5: data_out = 8'hBE;
                    16'hD9E6: data_out = 8'hBF;
                    16'hD9E7: data_out = 8'hC0;
                    16'hD9E8: data_out = 8'hC1;
                    16'hD9E9: data_out = 8'hC2;
                    16'hD9EA: data_out = 8'hC3;
                    16'hD9EB: data_out = 8'hC4;
                    16'hD9EC: data_out = 8'hC5;
                    16'hD9ED: data_out = 8'hC6;
                    16'hD9EE: data_out = 8'hC7;
                    16'hD9EF: data_out = 8'hC8;
                    16'hD9F0: data_out = 8'hC9;
                    16'hD9F1: data_out = 8'hCA;
                    16'hD9F2: data_out = 8'hCB;
                    16'hD9F3: data_out = 8'hCC;
                    16'hD9F4: data_out = 8'hCD;
                    16'hD9F5: data_out = 8'hCE;
                    16'hD9F6: data_out = 8'hCF;
                    16'hD9F7: data_out = 8'hD0;
                    16'hD9F8: data_out = 8'hD1;
                    16'hD9F9: data_out = 8'hD2;
                    16'hD9FA: data_out = 8'hD3;
                    16'hD9FB: data_out = 8'hD4;
                    16'hD9FC: data_out = 8'hD5;
                    16'hD9FD: data_out = 8'hD6;
                    16'hD9FE: data_out = 8'hD7;
                    16'hD9FF: data_out = 8'hD8;
                    16'hDA00: data_out = 8'hDA;
                    16'hDA01: data_out = 8'hD9;
                    16'hDA02: data_out = 8'hD8;
                    16'hDA03: data_out = 8'hD7;
                    16'hDA04: data_out = 8'hD6;
                    16'hDA05: data_out = 8'hD5;
                    16'hDA06: data_out = 8'hD4;
                    16'hDA07: data_out = 8'hD3;
                    16'hDA08: data_out = 8'hD2;
                    16'hDA09: data_out = 8'hD1;
                    16'hDA0A: data_out = 8'hD0;
                    16'hDA0B: data_out = 8'hCF;
                    16'hDA0C: data_out = 8'hCE;
                    16'hDA0D: data_out = 8'hCD;
                    16'hDA0E: data_out = 8'hCC;
                    16'hDA0F: data_out = 8'hCB;
                    16'hDA10: data_out = 8'hCA;
                    16'hDA11: data_out = 8'hC9;
                    16'hDA12: data_out = 8'hC8;
                    16'hDA13: data_out = 8'hC7;
                    16'hDA14: data_out = 8'hC6;
                    16'hDA15: data_out = 8'hC5;
                    16'hDA16: data_out = 8'hC4;
                    16'hDA17: data_out = 8'hC3;
                    16'hDA18: data_out = 8'hC2;
                    16'hDA19: data_out = 8'hC1;
                    16'hDA1A: data_out = 8'hC0;
                    16'hDA1B: data_out = 8'hBF;
                    16'hDA1C: data_out = 8'hBE;
                    16'hDA1D: data_out = 8'hBD;
                    16'hDA1E: data_out = 8'hBC;
                    16'hDA1F: data_out = 8'hBB;
                    16'hDA20: data_out = 8'hBA;
                    16'hDA21: data_out = 8'hB9;
                    16'hDA22: data_out = 8'hB8;
                    16'hDA23: data_out = 8'hB7;
                    16'hDA24: data_out = 8'hB6;
                    16'hDA25: data_out = 8'hB5;
                    16'hDA26: data_out = 8'hB4;
                    16'hDA27: data_out = 8'hB3;
                    16'hDA28: data_out = 8'hB2;
                    16'hDA29: data_out = 8'hB1;
                    16'hDA2A: data_out = 8'hB0;
                    16'hDA2B: data_out = 8'hAF;
                    16'hDA2C: data_out = 8'hAE;
                    16'hDA2D: data_out = 8'hAD;
                    16'hDA2E: data_out = 8'hAC;
                    16'hDA2F: data_out = 8'hAB;
                    16'hDA30: data_out = 8'hAA;
                    16'hDA31: data_out = 8'hA9;
                    16'hDA32: data_out = 8'hA8;
                    16'hDA33: data_out = 8'hA7;
                    16'hDA34: data_out = 8'hA6;
                    16'hDA35: data_out = 8'hA5;
                    16'hDA36: data_out = 8'hA4;
                    16'hDA37: data_out = 8'hA3;
                    16'hDA38: data_out = 8'hA2;
                    16'hDA39: data_out = 8'hA1;
                    16'hDA3A: data_out = 8'hA0;
                    16'hDA3B: data_out = 8'h9F;
                    16'hDA3C: data_out = 8'h9E;
                    16'hDA3D: data_out = 8'h9D;
                    16'hDA3E: data_out = 8'h9C;
                    16'hDA3F: data_out = 8'h9B;
                    16'hDA40: data_out = 8'h9A;
                    16'hDA41: data_out = 8'h99;
                    16'hDA42: data_out = 8'h98;
                    16'hDA43: data_out = 8'h97;
                    16'hDA44: data_out = 8'h96;
                    16'hDA45: data_out = 8'h95;
                    16'hDA46: data_out = 8'h94;
                    16'hDA47: data_out = 8'h93;
                    16'hDA48: data_out = 8'h92;
                    16'hDA49: data_out = 8'h91;
                    16'hDA4A: data_out = 8'h90;
                    16'hDA4B: data_out = 8'h8F;
                    16'hDA4C: data_out = 8'h8E;
                    16'hDA4D: data_out = 8'h8D;
                    16'hDA4E: data_out = 8'h8C;
                    16'hDA4F: data_out = 8'h8B;
                    16'hDA50: data_out = 8'h8A;
                    16'hDA51: data_out = 8'h89;
                    16'hDA52: data_out = 8'h88;
                    16'hDA53: data_out = 8'h87;
                    16'hDA54: data_out = 8'h86;
                    16'hDA55: data_out = 8'h85;
                    16'hDA56: data_out = 8'h84;
                    16'hDA57: data_out = 8'h83;
                    16'hDA58: data_out = 8'h82;
                    16'hDA59: data_out = 8'h81;
                    16'hDA5A: data_out = 8'h0;
                    16'hDA5B: data_out = 8'h1;
                    16'hDA5C: data_out = 8'h2;
                    16'hDA5D: data_out = 8'h3;
                    16'hDA5E: data_out = 8'h4;
                    16'hDA5F: data_out = 8'h5;
                    16'hDA60: data_out = 8'h6;
                    16'hDA61: data_out = 8'h7;
                    16'hDA62: data_out = 8'h8;
                    16'hDA63: data_out = 8'h9;
                    16'hDA64: data_out = 8'hA;
                    16'hDA65: data_out = 8'hB;
                    16'hDA66: data_out = 8'hC;
                    16'hDA67: data_out = 8'hD;
                    16'hDA68: data_out = 8'hE;
                    16'hDA69: data_out = 8'hF;
                    16'hDA6A: data_out = 8'h10;
                    16'hDA6B: data_out = 8'h11;
                    16'hDA6C: data_out = 8'h12;
                    16'hDA6D: data_out = 8'h13;
                    16'hDA6E: data_out = 8'h14;
                    16'hDA6F: data_out = 8'h15;
                    16'hDA70: data_out = 8'h16;
                    16'hDA71: data_out = 8'h17;
                    16'hDA72: data_out = 8'h18;
                    16'hDA73: data_out = 8'h19;
                    16'hDA74: data_out = 8'h1A;
                    16'hDA75: data_out = 8'h1B;
                    16'hDA76: data_out = 8'h1C;
                    16'hDA77: data_out = 8'h1D;
                    16'hDA78: data_out = 8'h1E;
                    16'hDA79: data_out = 8'h1F;
                    16'hDA7A: data_out = 8'h20;
                    16'hDA7B: data_out = 8'h21;
                    16'hDA7C: data_out = 8'h22;
                    16'hDA7D: data_out = 8'h23;
                    16'hDA7E: data_out = 8'h24;
                    16'hDA7F: data_out = 8'h25;
                    16'hDA80: data_out = 8'hDA;
                    16'hDA81: data_out = 8'hDB;
                    16'hDA82: data_out = 8'hDC;
                    16'hDA83: data_out = 8'hDD;
                    16'hDA84: data_out = 8'hDE;
                    16'hDA85: data_out = 8'hDF;
                    16'hDA86: data_out = 8'hE0;
                    16'hDA87: data_out = 8'hE1;
                    16'hDA88: data_out = 8'hE2;
                    16'hDA89: data_out = 8'hE3;
                    16'hDA8A: data_out = 8'hE4;
                    16'hDA8B: data_out = 8'hE5;
                    16'hDA8C: data_out = 8'hE6;
                    16'hDA8D: data_out = 8'hE7;
                    16'hDA8E: data_out = 8'hE8;
                    16'hDA8F: data_out = 8'hE9;
                    16'hDA90: data_out = 8'hEA;
                    16'hDA91: data_out = 8'hEB;
                    16'hDA92: data_out = 8'hEC;
                    16'hDA93: data_out = 8'hED;
                    16'hDA94: data_out = 8'hEE;
                    16'hDA95: data_out = 8'hEF;
                    16'hDA96: data_out = 8'hF0;
                    16'hDA97: data_out = 8'hF1;
                    16'hDA98: data_out = 8'hF2;
                    16'hDA99: data_out = 8'hF3;
                    16'hDA9A: data_out = 8'hF4;
                    16'hDA9B: data_out = 8'hF5;
                    16'hDA9C: data_out = 8'hF6;
                    16'hDA9D: data_out = 8'hF7;
                    16'hDA9E: data_out = 8'hF8;
                    16'hDA9F: data_out = 8'hF9;
                    16'hDAA0: data_out = 8'hFA;
                    16'hDAA1: data_out = 8'hFB;
                    16'hDAA2: data_out = 8'hFC;
                    16'hDAA3: data_out = 8'hFD;
                    16'hDAA4: data_out = 8'hFE;
                    16'hDAA5: data_out = 8'hFF;
                    16'hDAA6: data_out = 8'h80;
                    16'hDAA7: data_out = 8'h81;
                    16'hDAA8: data_out = 8'h82;
                    16'hDAA9: data_out = 8'h83;
                    16'hDAAA: data_out = 8'h84;
                    16'hDAAB: data_out = 8'h85;
                    16'hDAAC: data_out = 8'h86;
                    16'hDAAD: data_out = 8'h87;
                    16'hDAAE: data_out = 8'h88;
                    16'hDAAF: data_out = 8'h89;
                    16'hDAB0: data_out = 8'h8A;
                    16'hDAB1: data_out = 8'h8B;
                    16'hDAB2: data_out = 8'h8C;
                    16'hDAB3: data_out = 8'h8D;
                    16'hDAB4: data_out = 8'h8E;
                    16'hDAB5: data_out = 8'h8F;
                    16'hDAB6: data_out = 8'h90;
                    16'hDAB7: data_out = 8'h91;
                    16'hDAB8: data_out = 8'h92;
                    16'hDAB9: data_out = 8'h93;
                    16'hDABA: data_out = 8'h94;
                    16'hDABB: data_out = 8'h95;
                    16'hDABC: data_out = 8'h96;
                    16'hDABD: data_out = 8'h97;
                    16'hDABE: data_out = 8'h98;
                    16'hDABF: data_out = 8'h99;
                    16'hDAC0: data_out = 8'h9A;
                    16'hDAC1: data_out = 8'h9B;
                    16'hDAC2: data_out = 8'h9C;
                    16'hDAC3: data_out = 8'h9D;
                    16'hDAC4: data_out = 8'h9E;
                    16'hDAC5: data_out = 8'h9F;
                    16'hDAC6: data_out = 8'hA0;
                    16'hDAC7: data_out = 8'hA1;
                    16'hDAC8: data_out = 8'hA2;
                    16'hDAC9: data_out = 8'hA3;
                    16'hDACA: data_out = 8'hA4;
                    16'hDACB: data_out = 8'hA5;
                    16'hDACC: data_out = 8'hA6;
                    16'hDACD: data_out = 8'hA7;
                    16'hDACE: data_out = 8'hA8;
                    16'hDACF: data_out = 8'hA9;
                    16'hDAD0: data_out = 8'hAA;
                    16'hDAD1: data_out = 8'hAB;
                    16'hDAD2: data_out = 8'hAC;
                    16'hDAD3: data_out = 8'hAD;
                    16'hDAD4: data_out = 8'hAE;
                    16'hDAD5: data_out = 8'hAF;
                    16'hDAD6: data_out = 8'hB0;
                    16'hDAD7: data_out = 8'hB1;
                    16'hDAD8: data_out = 8'hB2;
                    16'hDAD9: data_out = 8'hB3;
                    16'hDADA: data_out = 8'hB4;
                    16'hDADB: data_out = 8'hB5;
                    16'hDADC: data_out = 8'hB6;
                    16'hDADD: data_out = 8'hB7;
                    16'hDADE: data_out = 8'hB8;
                    16'hDADF: data_out = 8'hB9;
                    16'hDAE0: data_out = 8'hBA;
                    16'hDAE1: data_out = 8'hBB;
                    16'hDAE2: data_out = 8'hBC;
                    16'hDAE3: data_out = 8'hBD;
                    16'hDAE4: data_out = 8'hBE;
                    16'hDAE5: data_out = 8'hBF;
                    16'hDAE6: data_out = 8'hC0;
                    16'hDAE7: data_out = 8'hC1;
                    16'hDAE8: data_out = 8'hC2;
                    16'hDAE9: data_out = 8'hC3;
                    16'hDAEA: data_out = 8'hC4;
                    16'hDAEB: data_out = 8'hC5;
                    16'hDAEC: data_out = 8'hC6;
                    16'hDAED: data_out = 8'hC7;
                    16'hDAEE: data_out = 8'hC8;
                    16'hDAEF: data_out = 8'hC9;
                    16'hDAF0: data_out = 8'hCA;
                    16'hDAF1: data_out = 8'hCB;
                    16'hDAF2: data_out = 8'hCC;
                    16'hDAF3: data_out = 8'hCD;
                    16'hDAF4: data_out = 8'hCE;
                    16'hDAF5: data_out = 8'hCF;
                    16'hDAF6: data_out = 8'hD0;
                    16'hDAF7: data_out = 8'hD1;
                    16'hDAF8: data_out = 8'hD2;
                    16'hDAF9: data_out = 8'hD3;
                    16'hDAFA: data_out = 8'hD4;
                    16'hDAFB: data_out = 8'hD5;
                    16'hDAFC: data_out = 8'hD6;
                    16'hDAFD: data_out = 8'hD7;
                    16'hDAFE: data_out = 8'hD8;
                    16'hDAFF: data_out = 8'hD9;
                    16'hDB00: data_out = 8'hDB;
                    16'hDB01: data_out = 8'hDA;
                    16'hDB02: data_out = 8'hD9;
                    16'hDB03: data_out = 8'hD8;
                    16'hDB04: data_out = 8'hD7;
                    16'hDB05: data_out = 8'hD6;
                    16'hDB06: data_out = 8'hD5;
                    16'hDB07: data_out = 8'hD4;
                    16'hDB08: data_out = 8'hD3;
                    16'hDB09: data_out = 8'hD2;
                    16'hDB0A: data_out = 8'hD1;
                    16'hDB0B: data_out = 8'hD0;
                    16'hDB0C: data_out = 8'hCF;
                    16'hDB0D: data_out = 8'hCE;
                    16'hDB0E: data_out = 8'hCD;
                    16'hDB0F: data_out = 8'hCC;
                    16'hDB10: data_out = 8'hCB;
                    16'hDB11: data_out = 8'hCA;
                    16'hDB12: data_out = 8'hC9;
                    16'hDB13: data_out = 8'hC8;
                    16'hDB14: data_out = 8'hC7;
                    16'hDB15: data_out = 8'hC6;
                    16'hDB16: data_out = 8'hC5;
                    16'hDB17: data_out = 8'hC4;
                    16'hDB18: data_out = 8'hC3;
                    16'hDB19: data_out = 8'hC2;
                    16'hDB1A: data_out = 8'hC1;
                    16'hDB1B: data_out = 8'hC0;
                    16'hDB1C: data_out = 8'hBF;
                    16'hDB1D: data_out = 8'hBE;
                    16'hDB1E: data_out = 8'hBD;
                    16'hDB1F: data_out = 8'hBC;
                    16'hDB20: data_out = 8'hBB;
                    16'hDB21: data_out = 8'hBA;
                    16'hDB22: data_out = 8'hB9;
                    16'hDB23: data_out = 8'hB8;
                    16'hDB24: data_out = 8'hB7;
                    16'hDB25: data_out = 8'hB6;
                    16'hDB26: data_out = 8'hB5;
                    16'hDB27: data_out = 8'hB4;
                    16'hDB28: data_out = 8'hB3;
                    16'hDB29: data_out = 8'hB2;
                    16'hDB2A: data_out = 8'hB1;
                    16'hDB2B: data_out = 8'hB0;
                    16'hDB2C: data_out = 8'hAF;
                    16'hDB2D: data_out = 8'hAE;
                    16'hDB2E: data_out = 8'hAD;
                    16'hDB2F: data_out = 8'hAC;
                    16'hDB30: data_out = 8'hAB;
                    16'hDB31: data_out = 8'hAA;
                    16'hDB32: data_out = 8'hA9;
                    16'hDB33: data_out = 8'hA8;
                    16'hDB34: data_out = 8'hA7;
                    16'hDB35: data_out = 8'hA6;
                    16'hDB36: data_out = 8'hA5;
                    16'hDB37: data_out = 8'hA4;
                    16'hDB38: data_out = 8'hA3;
                    16'hDB39: data_out = 8'hA2;
                    16'hDB3A: data_out = 8'hA1;
                    16'hDB3B: data_out = 8'hA0;
                    16'hDB3C: data_out = 8'h9F;
                    16'hDB3D: data_out = 8'h9E;
                    16'hDB3E: data_out = 8'h9D;
                    16'hDB3F: data_out = 8'h9C;
                    16'hDB40: data_out = 8'h9B;
                    16'hDB41: data_out = 8'h9A;
                    16'hDB42: data_out = 8'h99;
                    16'hDB43: data_out = 8'h98;
                    16'hDB44: data_out = 8'h97;
                    16'hDB45: data_out = 8'h96;
                    16'hDB46: data_out = 8'h95;
                    16'hDB47: data_out = 8'h94;
                    16'hDB48: data_out = 8'h93;
                    16'hDB49: data_out = 8'h92;
                    16'hDB4A: data_out = 8'h91;
                    16'hDB4B: data_out = 8'h90;
                    16'hDB4C: data_out = 8'h8F;
                    16'hDB4D: data_out = 8'h8E;
                    16'hDB4E: data_out = 8'h8D;
                    16'hDB4F: data_out = 8'h8C;
                    16'hDB50: data_out = 8'h8B;
                    16'hDB51: data_out = 8'h8A;
                    16'hDB52: data_out = 8'h89;
                    16'hDB53: data_out = 8'h88;
                    16'hDB54: data_out = 8'h87;
                    16'hDB55: data_out = 8'h86;
                    16'hDB56: data_out = 8'h85;
                    16'hDB57: data_out = 8'h84;
                    16'hDB58: data_out = 8'h83;
                    16'hDB59: data_out = 8'h82;
                    16'hDB5A: data_out = 8'h81;
                    16'hDB5B: data_out = 8'h0;
                    16'hDB5C: data_out = 8'h1;
                    16'hDB5D: data_out = 8'h2;
                    16'hDB5E: data_out = 8'h3;
                    16'hDB5F: data_out = 8'h4;
                    16'hDB60: data_out = 8'h5;
                    16'hDB61: data_out = 8'h6;
                    16'hDB62: data_out = 8'h7;
                    16'hDB63: data_out = 8'h8;
                    16'hDB64: data_out = 8'h9;
                    16'hDB65: data_out = 8'hA;
                    16'hDB66: data_out = 8'hB;
                    16'hDB67: data_out = 8'hC;
                    16'hDB68: data_out = 8'hD;
                    16'hDB69: data_out = 8'hE;
                    16'hDB6A: data_out = 8'hF;
                    16'hDB6B: data_out = 8'h10;
                    16'hDB6C: data_out = 8'h11;
                    16'hDB6D: data_out = 8'h12;
                    16'hDB6E: data_out = 8'h13;
                    16'hDB6F: data_out = 8'h14;
                    16'hDB70: data_out = 8'h15;
                    16'hDB71: data_out = 8'h16;
                    16'hDB72: data_out = 8'h17;
                    16'hDB73: data_out = 8'h18;
                    16'hDB74: data_out = 8'h19;
                    16'hDB75: data_out = 8'h1A;
                    16'hDB76: data_out = 8'h1B;
                    16'hDB77: data_out = 8'h1C;
                    16'hDB78: data_out = 8'h1D;
                    16'hDB79: data_out = 8'h1E;
                    16'hDB7A: data_out = 8'h1F;
                    16'hDB7B: data_out = 8'h20;
                    16'hDB7C: data_out = 8'h21;
                    16'hDB7D: data_out = 8'h22;
                    16'hDB7E: data_out = 8'h23;
                    16'hDB7F: data_out = 8'h24;
                    16'hDB80: data_out = 8'hDB;
                    16'hDB81: data_out = 8'hDC;
                    16'hDB82: data_out = 8'hDD;
                    16'hDB83: data_out = 8'hDE;
                    16'hDB84: data_out = 8'hDF;
                    16'hDB85: data_out = 8'hE0;
                    16'hDB86: data_out = 8'hE1;
                    16'hDB87: data_out = 8'hE2;
                    16'hDB88: data_out = 8'hE3;
                    16'hDB89: data_out = 8'hE4;
                    16'hDB8A: data_out = 8'hE5;
                    16'hDB8B: data_out = 8'hE6;
                    16'hDB8C: data_out = 8'hE7;
                    16'hDB8D: data_out = 8'hE8;
                    16'hDB8E: data_out = 8'hE9;
                    16'hDB8F: data_out = 8'hEA;
                    16'hDB90: data_out = 8'hEB;
                    16'hDB91: data_out = 8'hEC;
                    16'hDB92: data_out = 8'hED;
                    16'hDB93: data_out = 8'hEE;
                    16'hDB94: data_out = 8'hEF;
                    16'hDB95: data_out = 8'hF0;
                    16'hDB96: data_out = 8'hF1;
                    16'hDB97: data_out = 8'hF2;
                    16'hDB98: data_out = 8'hF3;
                    16'hDB99: data_out = 8'hF4;
                    16'hDB9A: data_out = 8'hF5;
                    16'hDB9B: data_out = 8'hF6;
                    16'hDB9C: data_out = 8'hF7;
                    16'hDB9D: data_out = 8'hF8;
                    16'hDB9E: data_out = 8'hF9;
                    16'hDB9F: data_out = 8'hFA;
                    16'hDBA0: data_out = 8'hFB;
                    16'hDBA1: data_out = 8'hFC;
                    16'hDBA2: data_out = 8'hFD;
                    16'hDBA3: data_out = 8'hFE;
                    16'hDBA4: data_out = 8'hFF;
                    16'hDBA5: data_out = 8'h80;
                    16'hDBA6: data_out = 8'h81;
                    16'hDBA7: data_out = 8'h82;
                    16'hDBA8: data_out = 8'h83;
                    16'hDBA9: data_out = 8'h84;
                    16'hDBAA: data_out = 8'h85;
                    16'hDBAB: data_out = 8'h86;
                    16'hDBAC: data_out = 8'h87;
                    16'hDBAD: data_out = 8'h88;
                    16'hDBAE: data_out = 8'h89;
                    16'hDBAF: data_out = 8'h8A;
                    16'hDBB0: data_out = 8'h8B;
                    16'hDBB1: data_out = 8'h8C;
                    16'hDBB2: data_out = 8'h8D;
                    16'hDBB3: data_out = 8'h8E;
                    16'hDBB4: data_out = 8'h8F;
                    16'hDBB5: data_out = 8'h90;
                    16'hDBB6: data_out = 8'h91;
                    16'hDBB7: data_out = 8'h92;
                    16'hDBB8: data_out = 8'h93;
                    16'hDBB9: data_out = 8'h94;
                    16'hDBBA: data_out = 8'h95;
                    16'hDBBB: data_out = 8'h96;
                    16'hDBBC: data_out = 8'h97;
                    16'hDBBD: data_out = 8'h98;
                    16'hDBBE: data_out = 8'h99;
                    16'hDBBF: data_out = 8'h9A;
                    16'hDBC0: data_out = 8'h9B;
                    16'hDBC1: data_out = 8'h9C;
                    16'hDBC2: data_out = 8'h9D;
                    16'hDBC3: data_out = 8'h9E;
                    16'hDBC4: data_out = 8'h9F;
                    16'hDBC5: data_out = 8'hA0;
                    16'hDBC6: data_out = 8'hA1;
                    16'hDBC7: data_out = 8'hA2;
                    16'hDBC8: data_out = 8'hA3;
                    16'hDBC9: data_out = 8'hA4;
                    16'hDBCA: data_out = 8'hA5;
                    16'hDBCB: data_out = 8'hA6;
                    16'hDBCC: data_out = 8'hA7;
                    16'hDBCD: data_out = 8'hA8;
                    16'hDBCE: data_out = 8'hA9;
                    16'hDBCF: data_out = 8'hAA;
                    16'hDBD0: data_out = 8'hAB;
                    16'hDBD1: data_out = 8'hAC;
                    16'hDBD2: data_out = 8'hAD;
                    16'hDBD3: data_out = 8'hAE;
                    16'hDBD4: data_out = 8'hAF;
                    16'hDBD5: data_out = 8'hB0;
                    16'hDBD6: data_out = 8'hB1;
                    16'hDBD7: data_out = 8'hB2;
                    16'hDBD8: data_out = 8'hB3;
                    16'hDBD9: data_out = 8'hB4;
                    16'hDBDA: data_out = 8'hB5;
                    16'hDBDB: data_out = 8'hB6;
                    16'hDBDC: data_out = 8'hB7;
                    16'hDBDD: data_out = 8'hB8;
                    16'hDBDE: data_out = 8'hB9;
                    16'hDBDF: data_out = 8'hBA;
                    16'hDBE0: data_out = 8'hBB;
                    16'hDBE1: data_out = 8'hBC;
                    16'hDBE2: data_out = 8'hBD;
                    16'hDBE3: data_out = 8'hBE;
                    16'hDBE4: data_out = 8'hBF;
                    16'hDBE5: data_out = 8'hC0;
                    16'hDBE6: data_out = 8'hC1;
                    16'hDBE7: data_out = 8'hC2;
                    16'hDBE8: data_out = 8'hC3;
                    16'hDBE9: data_out = 8'hC4;
                    16'hDBEA: data_out = 8'hC5;
                    16'hDBEB: data_out = 8'hC6;
                    16'hDBEC: data_out = 8'hC7;
                    16'hDBED: data_out = 8'hC8;
                    16'hDBEE: data_out = 8'hC9;
                    16'hDBEF: data_out = 8'hCA;
                    16'hDBF0: data_out = 8'hCB;
                    16'hDBF1: data_out = 8'hCC;
                    16'hDBF2: data_out = 8'hCD;
                    16'hDBF3: data_out = 8'hCE;
                    16'hDBF4: data_out = 8'hCF;
                    16'hDBF5: data_out = 8'hD0;
                    16'hDBF6: data_out = 8'hD1;
                    16'hDBF7: data_out = 8'hD2;
                    16'hDBF8: data_out = 8'hD3;
                    16'hDBF9: data_out = 8'hD4;
                    16'hDBFA: data_out = 8'hD5;
                    16'hDBFB: data_out = 8'hD6;
                    16'hDBFC: data_out = 8'hD7;
                    16'hDBFD: data_out = 8'hD8;
                    16'hDBFE: data_out = 8'hD9;
                    16'hDBFF: data_out = 8'hDA;
                    16'hDC00: data_out = 8'hDC;
                    16'hDC01: data_out = 8'hDB;
                    16'hDC02: data_out = 8'hDA;
                    16'hDC03: data_out = 8'hD9;
                    16'hDC04: data_out = 8'hD8;
                    16'hDC05: data_out = 8'hD7;
                    16'hDC06: data_out = 8'hD6;
                    16'hDC07: data_out = 8'hD5;
                    16'hDC08: data_out = 8'hD4;
                    16'hDC09: data_out = 8'hD3;
                    16'hDC0A: data_out = 8'hD2;
                    16'hDC0B: data_out = 8'hD1;
                    16'hDC0C: data_out = 8'hD0;
                    16'hDC0D: data_out = 8'hCF;
                    16'hDC0E: data_out = 8'hCE;
                    16'hDC0F: data_out = 8'hCD;
                    16'hDC10: data_out = 8'hCC;
                    16'hDC11: data_out = 8'hCB;
                    16'hDC12: data_out = 8'hCA;
                    16'hDC13: data_out = 8'hC9;
                    16'hDC14: data_out = 8'hC8;
                    16'hDC15: data_out = 8'hC7;
                    16'hDC16: data_out = 8'hC6;
                    16'hDC17: data_out = 8'hC5;
                    16'hDC18: data_out = 8'hC4;
                    16'hDC19: data_out = 8'hC3;
                    16'hDC1A: data_out = 8'hC2;
                    16'hDC1B: data_out = 8'hC1;
                    16'hDC1C: data_out = 8'hC0;
                    16'hDC1D: data_out = 8'hBF;
                    16'hDC1E: data_out = 8'hBE;
                    16'hDC1F: data_out = 8'hBD;
                    16'hDC20: data_out = 8'hBC;
                    16'hDC21: data_out = 8'hBB;
                    16'hDC22: data_out = 8'hBA;
                    16'hDC23: data_out = 8'hB9;
                    16'hDC24: data_out = 8'hB8;
                    16'hDC25: data_out = 8'hB7;
                    16'hDC26: data_out = 8'hB6;
                    16'hDC27: data_out = 8'hB5;
                    16'hDC28: data_out = 8'hB4;
                    16'hDC29: data_out = 8'hB3;
                    16'hDC2A: data_out = 8'hB2;
                    16'hDC2B: data_out = 8'hB1;
                    16'hDC2C: data_out = 8'hB0;
                    16'hDC2D: data_out = 8'hAF;
                    16'hDC2E: data_out = 8'hAE;
                    16'hDC2F: data_out = 8'hAD;
                    16'hDC30: data_out = 8'hAC;
                    16'hDC31: data_out = 8'hAB;
                    16'hDC32: data_out = 8'hAA;
                    16'hDC33: data_out = 8'hA9;
                    16'hDC34: data_out = 8'hA8;
                    16'hDC35: data_out = 8'hA7;
                    16'hDC36: data_out = 8'hA6;
                    16'hDC37: data_out = 8'hA5;
                    16'hDC38: data_out = 8'hA4;
                    16'hDC39: data_out = 8'hA3;
                    16'hDC3A: data_out = 8'hA2;
                    16'hDC3B: data_out = 8'hA1;
                    16'hDC3C: data_out = 8'hA0;
                    16'hDC3D: data_out = 8'h9F;
                    16'hDC3E: data_out = 8'h9E;
                    16'hDC3F: data_out = 8'h9D;
                    16'hDC40: data_out = 8'h9C;
                    16'hDC41: data_out = 8'h9B;
                    16'hDC42: data_out = 8'h9A;
                    16'hDC43: data_out = 8'h99;
                    16'hDC44: data_out = 8'h98;
                    16'hDC45: data_out = 8'h97;
                    16'hDC46: data_out = 8'h96;
                    16'hDC47: data_out = 8'h95;
                    16'hDC48: data_out = 8'h94;
                    16'hDC49: data_out = 8'h93;
                    16'hDC4A: data_out = 8'h92;
                    16'hDC4B: data_out = 8'h91;
                    16'hDC4C: data_out = 8'h90;
                    16'hDC4D: data_out = 8'h8F;
                    16'hDC4E: data_out = 8'h8E;
                    16'hDC4F: data_out = 8'h8D;
                    16'hDC50: data_out = 8'h8C;
                    16'hDC51: data_out = 8'h8B;
                    16'hDC52: data_out = 8'h8A;
                    16'hDC53: data_out = 8'h89;
                    16'hDC54: data_out = 8'h88;
                    16'hDC55: data_out = 8'h87;
                    16'hDC56: data_out = 8'h86;
                    16'hDC57: data_out = 8'h85;
                    16'hDC58: data_out = 8'h84;
                    16'hDC59: data_out = 8'h83;
                    16'hDC5A: data_out = 8'h82;
                    16'hDC5B: data_out = 8'h81;
                    16'hDC5C: data_out = 8'h0;
                    16'hDC5D: data_out = 8'h1;
                    16'hDC5E: data_out = 8'h2;
                    16'hDC5F: data_out = 8'h3;
                    16'hDC60: data_out = 8'h4;
                    16'hDC61: data_out = 8'h5;
                    16'hDC62: data_out = 8'h6;
                    16'hDC63: data_out = 8'h7;
                    16'hDC64: data_out = 8'h8;
                    16'hDC65: data_out = 8'h9;
                    16'hDC66: data_out = 8'hA;
                    16'hDC67: data_out = 8'hB;
                    16'hDC68: data_out = 8'hC;
                    16'hDC69: data_out = 8'hD;
                    16'hDC6A: data_out = 8'hE;
                    16'hDC6B: data_out = 8'hF;
                    16'hDC6C: data_out = 8'h10;
                    16'hDC6D: data_out = 8'h11;
                    16'hDC6E: data_out = 8'h12;
                    16'hDC6F: data_out = 8'h13;
                    16'hDC70: data_out = 8'h14;
                    16'hDC71: data_out = 8'h15;
                    16'hDC72: data_out = 8'h16;
                    16'hDC73: data_out = 8'h17;
                    16'hDC74: data_out = 8'h18;
                    16'hDC75: data_out = 8'h19;
                    16'hDC76: data_out = 8'h1A;
                    16'hDC77: data_out = 8'h1B;
                    16'hDC78: data_out = 8'h1C;
                    16'hDC79: data_out = 8'h1D;
                    16'hDC7A: data_out = 8'h1E;
                    16'hDC7B: data_out = 8'h1F;
                    16'hDC7C: data_out = 8'h20;
                    16'hDC7D: data_out = 8'h21;
                    16'hDC7E: data_out = 8'h22;
                    16'hDC7F: data_out = 8'h23;
                    16'hDC80: data_out = 8'hDC;
                    16'hDC81: data_out = 8'hDD;
                    16'hDC82: data_out = 8'hDE;
                    16'hDC83: data_out = 8'hDF;
                    16'hDC84: data_out = 8'hE0;
                    16'hDC85: data_out = 8'hE1;
                    16'hDC86: data_out = 8'hE2;
                    16'hDC87: data_out = 8'hE3;
                    16'hDC88: data_out = 8'hE4;
                    16'hDC89: data_out = 8'hE5;
                    16'hDC8A: data_out = 8'hE6;
                    16'hDC8B: data_out = 8'hE7;
                    16'hDC8C: data_out = 8'hE8;
                    16'hDC8D: data_out = 8'hE9;
                    16'hDC8E: data_out = 8'hEA;
                    16'hDC8F: data_out = 8'hEB;
                    16'hDC90: data_out = 8'hEC;
                    16'hDC91: data_out = 8'hED;
                    16'hDC92: data_out = 8'hEE;
                    16'hDC93: data_out = 8'hEF;
                    16'hDC94: data_out = 8'hF0;
                    16'hDC95: data_out = 8'hF1;
                    16'hDC96: data_out = 8'hF2;
                    16'hDC97: data_out = 8'hF3;
                    16'hDC98: data_out = 8'hF4;
                    16'hDC99: data_out = 8'hF5;
                    16'hDC9A: data_out = 8'hF6;
                    16'hDC9B: data_out = 8'hF7;
                    16'hDC9C: data_out = 8'hF8;
                    16'hDC9D: data_out = 8'hF9;
                    16'hDC9E: data_out = 8'hFA;
                    16'hDC9F: data_out = 8'hFB;
                    16'hDCA0: data_out = 8'hFC;
                    16'hDCA1: data_out = 8'hFD;
                    16'hDCA2: data_out = 8'hFE;
                    16'hDCA3: data_out = 8'hFF;
                    16'hDCA4: data_out = 8'h80;
                    16'hDCA5: data_out = 8'h81;
                    16'hDCA6: data_out = 8'h82;
                    16'hDCA7: data_out = 8'h83;
                    16'hDCA8: data_out = 8'h84;
                    16'hDCA9: data_out = 8'h85;
                    16'hDCAA: data_out = 8'h86;
                    16'hDCAB: data_out = 8'h87;
                    16'hDCAC: data_out = 8'h88;
                    16'hDCAD: data_out = 8'h89;
                    16'hDCAE: data_out = 8'h8A;
                    16'hDCAF: data_out = 8'h8B;
                    16'hDCB0: data_out = 8'h8C;
                    16'hDCB1: data_out = 8'h8D;
                    16'hDCB2: data_out = 8'h8E;
                    16'hDCB3: data_out = 8'h8F;
                    16'hDCB4: data_out = 8'h90;
                    16'hDCB5: data_out = 8'h91;
                    16'hDCB6: data_out = 8'h92;
                    16'hDCB7: data_out = 8'h93;
                    16'hDCB8: data_out = 8'h94;
                    16'hDCB9: data_out = 8'h95;
                    16'hDCBA: data_out = 8'h96;
                    16'hDCBB: data_out = 8'h97;
                    16'hDCBC: data_out = 8'h98;
                    16'hDCBD: data_out = 8'h99;
                    16'hDCBE: data_out = 8'h9A;
                    16'hDCBF: data_out = 8'h9B;
                    16'hDCC0: data_out = 8'h9C;
                    16'hDCC1: data_out = 8'h9D;
                    16'hDCC2: data_out = 8'h9E;
                    16'hDCC3: data_out = 8'h9F;
                    16'hDCC4: data_out = 8'hA0;
                    16'hDCC5: data_out = 8'hA1;
                    16'hDCC6: data_out = 8'hA2;
                    16'hDCC7: data_out = 8'hA3;
                    16'hDCC8: data_out = 8'hA4;
                    16'hDCC9: data_out = 8'hA5;
                    16'hDCCA: data_out = 8'hA6;
                    16'hDCCB: data_out = 8'hA7;
                    16'hDCCC: data_out = 8'hA8;
                    16'hDCCD: data_out = 8'hA9;
                    16'hDCCE: data_out = 8'hAA;
                    16'hDCCF: data_out = 8'hAB;
                    16'hDCD0: data_out = 8'hAC;
                    16'hDCD1: data_out = 8'hAD;
                    16'hDCD2: data_out = 8'hAE;
                    16'hDCD3: data_out = 8'hAF;
                    16'hDCD4: data_out = 8'hB0;
                    16'hDCD5: data_out = 8'hB1;
                    16'hDCD6: data_out = 8'hB2;
                    16'hDCD7: data_out = 8'hB3;
                    16'hDCD8: data_out = 8'hB4;
                    16'hDCD9: data_out = 8'hB5;
                    16'hDCDA: data_out = 8'hB6;
                    16'hDCDB: data_out = 8'hB7;
                    16'hDCDC: data_out = 8'hB8;
                    16'hDCDD: data_out = 8'hB9;
                    16'hDCDE: data_out = 8'hBA;
                    16'hDCDF: data_out = 8'hBB;
                    16'hDCE0: data_out = 8'hBC;
                    16'hDCE1: data_out = 8'hBD;
                    16'hDCE2: data_out = 8'hBE;
                    16'hDCE3: data_out = 8'hBF;
                    16'hDCE4: data_out = 8'hC0;
                    16'hDCE5: data_out = 8'hC1;
                    16'hDCE6: data_out = 8'hC2;
                    16'hDCE7: data_out = 8'hC3;
                    16'hDCE8: data_out = 8'hC4;
                    16'hDCE9: data_out = 8'hC5;
                    16'hDCEA: data_out = 8'hC6;
                    16'hDCEB: data_out = 8'hC7;
                    16'hDCEC: data_out = 8'hC8;
                    16'hDCED: data_out = 8'hC9;
                    16'hDCEE: data_out = 8'hCA;
                    16'hDCEF: data_out = 8'hCB;
                    16'hDCF0: data_out = 8'hCC;
                    16'hDCF1: data_out = 8'hCD;
                    16'hDCF2: data_out = 8'hCE;
                    16'hDCF3: data_out = 8'hCF;
                    16'hDCF4: data_out = 8'hD0;
                    16'hDCF5: data_out = 8'hD1;
                    16'hDCF6: data_out = 8'hD2;
                    16'hDCF7: data_out = 8'hD3;
                    16'hDCF8: data_out = 8'hD4;
                    16'hDCF9: data_out = 8'hD5;
                    16'hDCFA: data_out = 8'hD6;
                    16'hDCFB: data_out = 8'hD7;
                    16'hDCFC: data_out = 8'hD8;
                    16'hDCFD: data_out = 8'hD9;
                    16'hDCFE: data_out = 8'hDA;
                    16'hDCFF: data_out = 8'hDB;
                    16'hDD00: data_out = 8'hDD;
                    16'hDD01: data_out = 8'hDC;
                    16'hDD02: data_out = 8'hDB;
                    16'hDD03: data_out = 8'hDA;
                    16'hDD04: data_out = 8'hD9;
                    16'hDD05: data_out = 8'hD8;
                    16'hDD06: data_out = 8'hD7;
                    16'hDD07: data_out = 8'hD6;
                    16'hDD08: data_out = 8'hD5;
                    16'hDD09: data_out = 8'hD4;
                    16'hDD0A: data_out = 8'hD3;
                    16'hDD0B: data_out = 8'hD2;
                    16'hDD0C: data_out = 8'hD1;
                    16'hDD0D: data_out = 8'hD0;
                    16'hDD0E: data_out = 8'hCF;
                    16'hDD0F: data_out = 8'hCE;
                    16'hDD10: data_out = 8'hCD;
                    16'hDD11: data_out = 8'hCC;
                    16'hDD12: data_out = 8'hCB;
                    16'hDD13: data_out = 8'hCA;
                    16'hDD14: data_out = 8'hC9;
                    16'hDD15: data_out = 8'hC8;
                    16'hDD16: data_out = 8'hC7;
                    16'hDD17: data_out = 8'hC6;
                    16'hDD18: data_out = 8'hC5;
                    16'hDD19: data_out = 8'hC4;
                    16'hDD1A: data_out = 8'hC3;
                    16'hDD1B: data_out = 8'hC2;
                    16'hDD1C: data_out = 8'hC1;
                    16'hDD1D: data_out = 8'hC0;
                    16'hDD1E: data_out = 8'hBF;
                    16'hDD1F: data_out = 8'hBE;
                    16'hDD20: data_out = 8'hBD;
                    16'hDD21: data_out = 8'hBC;
                    16'hDD22: data_out = 8'hBB;
                    16'hDD23: data_out = 8'hBA;
                    16'hDD24: data_out = 8'hB9;
                    16'hDD25: data_out = 8'hB8;
                    16'hDD26: data_out = 8'hB7;
                    16'hDD27: data_out = 8'hB6;
                    16'hDD28: data_out = 8'hB5;
                    16'hDD29: data_out = 8'hB4;
                    16'hDD2A: data_out = 8'hB3;
                    16'hDD2B: data_out = 8'hB2;
                    16'hDD2C: data_out = 8'hB1;
                    16'hDD2D: data_out = 8'hB0;
                    16'hDD2E: data_out = 8'hAF;
                    16'hDD2F: data_out = 8'hAE;
                    16'hDD30: data_out = 8'hAD;
                    16'hDD31: data_out = 8'hAC;
                    16'hDD32: data_out = 8'hAB;
                    16'hDD33: data_out = 8'hAA;
                    16'hDD34: data_out = 8'hA9;
                    16'hDD35: data_out = 8'hA8;
                    16'hDD36: data_out = 8'hA7;
                    16'hDD37: data_out = 8'hA6;
                    16'hDD38: data_out = 8'hA5;
                    16'hDD39: data_out = 8'hA4;
                    16'hDD3A: data_out = 8'hA3;
                    16'hDD3B: data_out = 8'hA2;
                    16'hDD3C: data_out = 8'hA1;
                    16'hDD3D: data_out = 8'hA0;
                    16'hDD3E: data_out = 8'h9F;
                    16'hDD3F: data_out = 8'h9E;
                    16'hDD40: data_out = 8'h9D;
                    16'hDD41: data_out = 8'h9C;
                    16'hDD42: data_out = 8'h9B;
                    16'hDD43: data_out = 8'h9A;
                    16'hDD44: data_out = 8'h99;
                    16'hDD45: data_out = 8'h98;
                    16'hDD46: data_out = 8'h97;
                    16'hDD47: data_out = 8'h96;
                    16'hDD48: data_out = 8'h95;
                    16'hDD49: data_out = 8'h94;
                    16'hDD4A: data_out = 8'h93;
                    16'hDD4B: data_out = 8'h92;
                    16'hDD4C: data_out = 8'h91;
                    16'hDD4D: data_out = 8'h90;
                    16'hDD4E: data_out = 8'h8F;
                    16'hDD4F: data_out = 8'h8E;
                    16'hDD50: data_out = 8'h8D;
                    16'hDD51: data_out = 8'h8C;
                    16'hDD52: data_out = 8'h8B;
                    16'hDD53: data_out = 8'h8A;
                    16'hDD54: data_out = 8'h89;
                    16'hDD55: data_out = 8'h88;
                    16'hDD56: data_out = 8'h87;
                    16'hDD57: data_out = 8'h86;
                    16'hDD58: data_out = 8'h85;
                    16'hDD59: data_out = 8'h84;
                    16'hDD5A: data_out = 8'h83;
                    16'hDD5B: data_out = 8'h82;
                    16'hDD5C: data_out = 8'h81;
                    16'hDD5D: data_out = 8'h0;
                    16'hDD5E: data_out = 8'h1;
                    16'hDD5F: data_out = 8'h2;
                    16'hDD60: data_out = 8'h3;
                    16'hDD61: data_out = 8'h4;
                    16'hDD62: data_out = 8'h5;
                    16'hDD63: data_out = 8'h6;
                    16'hDD64: data_out = 8'h7;
                    16'hDD65: data_out = 8'h8;
                    16'hDD66: data_out = 8'h9;
                    16'hDD67: data_out = 8'hA;
                    16'hDD68: data_out = 8'hB;
                    16'hDD69: data_out = 8'hC;
                    16'hDD6A: data_out = 8'hD;
                    16'hDD6B: data_out = 8'hE;
                    16'hDD6C: data_out = 8'hF;
                    16'hDD6D: data_out = 8'h10;
                    16'hDD6E: data_out = 8'h11;
                    16'hDD6F: data_out = 8'h12;
                    16'hDD70: data_out = 8'h13;
                    16'hDD71: data_out = 8'h14;
                    16'hDD72: data_out = 8'h15;
                    16'hDD73: data_out = 8'h16;
                    16'hDD74: data_out = 8'h17;
                    16'hDD75: data_out = 8'h18;
                    16'hDD76: data_out = 8'h19;
                    16'hDD77: data_out = 8'h1A;
                    16'hDD78: data_out = 8'h1B;
                    16'hDD79: data_out = 8'h1C;
                    16'hDD7A: data_out = 8'h1D;
                    16'hDD7B: data_out = 8'h1E;
                    16'hDD7C: data_out = 8'h1F;
                    16'hDD7D: data_out = 8'h20;
                    16'hDD7E: data_out = 8'h21;
                    16'hDD7F: data_out = 8'h22;
                    16'hDD80: data_out = 8'hDD;
                    16'hDD81: data_out = 8'hDE;
                    16'hDD82: data_out = 8'hDF;
                    16'hDD83: data_out = 8'hE0;
                    16'hDD84: data_out = 8'hE1;
                    16'hDD85: data_out = 8'hE2;
                    16'hDD86: data_out = 8'hE3;
                    16'hDD87: data_out = 8'hE4;
                    16'hDD88: data_out = 8'hE5;
                    16'hDD89: data_out = 8'hE6;
                    16'hDD8A: data_out = 8'hE7;
                    16'hDD8B: data_out = 8'hE8;
                    16'hDD8C: data_out = 8'hE9;
                    16'hDD8D: data_out = 8'hEA;
                    16'hDD8E: data_out = 8'hEB;
                    16'hDD8F: data_out = 8'hEC;
                    16'hDD90: data_out = 8'hED;
                    16'hDD91: data_out = 8'hEE;
                    16'hDD92: data_out = 8'hEF;
                    16'hDD93: data_out = 8'hF0;
                    16'hDD94: data_out = 8'hF1;
                    16'hDD95: data_out = 8'hF2;
                    16'hDD96: data_out = 8'hF3;
                    16'hDD97: data_out = 8'hF4;
                    16'hDD98: data_out = 8'hF5;
                    16'hDD99: data_out = 8'hF6;
                    16'hDD9A: data_out = 8'hF7;
                    16'hDD9B: data_out = 8'hF8;
                    16'hDD9C: data_out = 8'hF9;
                    16'hDD9D: data_out = 8'hFA;
                    16'hDD9E: data_out = 8'hFB;
                    16'hDD9F: data_out = 8'hFC;
                    16'hDDA0: data_out = 8'hFD;
                    16'hDDA1: data_out = 8'hFE;
                    16'hDDA2: data_out = 8'hFF;
                    16'hDDA3: data_out = 8'h80;
                    16'hDDA4: data_out = 8'h81;
                    16'hDDA5: data_out = 8'h82;
                    16'hDDA6: data_out = 8'h83;
                    16'hDDA7: data_out = 8'h84;
                    16'hDDA8: data_out = 8'h85;
                    16'hDDA9: data_out = 8'h86;
                    16'hDDAA: data_out = 8'h87;
                    16'hDDAB: data_out = 8'h88;
                    16'hDDAC: data_out = 8'h89;
                    16'hDDAD: data_out = 8'h8A;
                    16'hDDAE: data_out = 8'h8B;
                    16'hDDAF: data_out = 8'h8C;
                    16'hDDB0: data_out = 8'h8D;
                    16'hDDB1: data_out = 8'h8E;
                    16'hDDB2: data_out = 8'h8F;
                    16'hDDB3: data_out = 8'h90;
                    16'hDDB4: data_out = 8'h91;
                    16'hDDB5: data_out = 8'h92;
                    16'hDDB6: data_out = 8'h93;
                    16'hDDB7: data_out = 8'h94;
                    16'hDDB8: data_out = 8'h95;
                    16'hDDB9: data_out = 8'h96;
                    16'hDDBA: data_out = 8'h97;
                    16'hDDBB: data_out = 8'h98;
                    16'hDDBC: data_out = 8'h99;
                    16'hDDBD: data_out = 8'h9A;
                    16'hDDBE: data_out = 8'h9B;
                    16'hDDBF: data_out = 8'h9C;
                    16'hDDC0: data_out = 8'h9D;
                    16'hDDC1: data_out = 8'h9E;
                    16'hDDC2: data_out = 8'h9F;
                    16'hDDC3: data_out = 8'hA0;
                    16'hDDC4: data_out = 8'hA1;
                    16'hDDC5: data_out = 8'hA2;
                    16'hDDC6: data_out = 8'hA3;
                    16'hDDC7: data_out = 8'hA4;
                    16'hDDC8: data_out = 8'hA5;
                    16'hDDC9: data_out = 8'hA6;
                    16'hDDCA: data_out = 8'hA7;
                    16'hDDCB: data_out = 8'hA8;
                    16'hDDCC: data_out = 8'hA9;
                    16'hDDCD: data_out = 8'hAA;
                    16'hDDCE: data_out = 8'hAB;
                    16'hDDCF: data_out = 8'hAC;
                    16'hDDD0: data_out = 8'hAD;
                    16'hDDD1: data_out = 8'hAE;
                    16'hDDD2: data_out = 8'hAF;
                    16'hDDD3: data_out = 8'hB0;
                    16'hDDD4: data_out = 8'hB1;
                    16'hDDD5: data_out = 8'hB2;
                    16'hDDD6: data_out = 8'hB3;
                    16'hDDD7: data_out = 8'hB4;
                    16'hDDD8: data_out = 8'hB5;
                    16'hDDD9: data_out = 8'hB6;
                    16'hDDDA: data_out = 8'hB7;
                    16'hDDDB: data_out = 8'hB8;
                    16'hDDDC: data_out = 8'hB9;
                    16'hDDDD: data_out = 8'hBA;
                    16'hDDDE: data_out = 8'hBB;
                    16'hDDDF: data_out = 8'hBC;
                    16'hDDE0: data_out = 8'hBD;
                    16'hDDE1: data_out = 8'hBE;
                    16'hDDE2: data_out = 8'hBF;
                    16'hDDE3: data_out = 8'hC0;
                    16'hDDE4: data_out = 8'hC1;
                    16'hDDE5: data_out = 8'hC2;
                    16'hDDE6: data_out = 8'hC3;
                    16'hDDE7: data_out = 8'hC4;
                    16'hDDE8: data_out = 8'hC5;
                    16'hDDE9: data_out = 8'hC6;
                    16'hDDEA: data_out = 8'hC7;
                    16'hDDEB: data_out = 8'hC8;
                    16'hDDEC: data_out = 8'hC9;
                    16'hDDED: data_out = 8'hCA;
                    16'hDDEE: data_out = 8'hCB;
                    16'hDDEF: data_out = 8'hCC;
                    16'hDDF0: data_out = 8'hCD;
                    16'hDDF1: data_out = 8'hCE;
                    16'hDDF2: data_out = 8'hCF;
                    16'hDDF3: data_out = 8'hD0;
                    16'hDDF4: data_out = 8'hD1;
                    16'hDDF5: data_out = 8'hD2;
                    16'hDDF6: data_out = 8'hD3;
                    16'hDDF7: data_out = 8'hD4;
                    16'hDDF8: data_out = 8'hD5;
                    16'hDDF9: data_out = 8'hD6;
                    16'hDDFA: data_out = 8'hD7;
                    16'hDDFB: data_out = 8'hD8;
                    16'hDDFC: data_out = 8'hD9;
                    16'hDDFD: data_out = 8'hDA;
                    16'hDDFE: data_out = 8'hDB;
                    16'hDDFF: data_out = 8'hDC;
                    16'hDE00: data_out = 8'hDE;
                    16'hDE01: data_out = 8'hDD;
                    16'hDE02: data_out = 8'hDC;
                    16'hDE03: data_out = 8'hDB;
                    16'hDE04: data_out = 8'hDA;
                    16'hDE05: data_out = 8'hD9;
                    16'hDE06: data_out = 8'hD8;
                    16'hDE07: data_out = 8'hD7;
                    16'hDE08: data_out = 8'hD6;
                    16'hDE09: data_out = 8'hD5;
                    16'hDE0A: data_out = 8'hD4;
                    16'hDE0B: data_out = 8'hD3;
                    16'hDE0C: data_out = 8'hD2;
                    16'hDE0D: data_out = 8'hD1;
                    16'hDE0E: data_out = 8'hD0;
                    16'hDE0F: data_out = 8'hCF;
                    16'hDE10: data_out = 8'hCE;
                    16'hDE11: data_out = 8'hCD;
                    16'hDE12: data_out = 8'hCC;
                    16'hDE13: data_out = 8'hCB;
                    16'hDE14: data_out = 8'hCA;
                    16'hDE15: data_out = 8'hC9;
                    16'hDE16: data_out = 8'hC8;
                    16'hDE17: data_out = 8'hC7;
                    16'hDE18: data_out = 8'hC6;
                    16'hDE19: data_out = 8'hC5;
                    16'hDE1A: data_out = 8'hC4;
                    16'hDE1B: data_out = 8'hC3;
                    16'hDE1C: data_out = 8'hC2;
                    16'hDE1D: data_out = 8'hC1;
                    16'hDE1E: data_out = 8'hC0;
                    16'hDE1F: data_out = 8'hBF;
                    16'hDE20: data_out = 8'hBE;
                    16'hDE21: data_out = 8'hBD;
                    16'hDE22: data_out = 8'hBC;
                    16'hDE23: data_out = 8'hBB;
                    16'hDE24: data_out = 8'hBA;
                    16'hDE25: data_out = 8'hB9;
                    16'hDE26: data_out = 8'hB8;
                    16'hDE27: data_out = 8'hB7;
                    16'hDE28: data_out = 8'hB6;
                    16'hDE29: data_out = 8'hB5;
                    16'hDE2A: data_out = 8'hB4;
                    16'hDE2B: data_out = 8'hB3;
                    16'hDE2C: data_out = 8'hB2;
                    16'hDE2D: data_out = 8'hB1;
                    16'hDE2E: data_out = 8'hB0;
                    16'hDE2F: data_out = 8'hAF;
                    16'hDE30: data_out = 8'hAE;
                    16'hDE31: data_out = 8'hAD;
                    16'hDE32: data_out = 8'hAC;
                    16'hDE33: data_out = 8'hAB;
                    16'hDE34: data_out = 8'hAA;
                    16'hDE35: data_out = 8'hA9;
                    16'hDE36: data_out = 8'hA8;
                    16'hDE37: data_out = 8'hA7;
                    16'hDE38: data_out = 8'hA6;
                    16'hDE39: data_out = 8'hA5;
                    16'hDE3A: data_out = 8'hA4;
                    16'hDE3B: data_out = 8'hA3;
                    16'hDE3C: data_out = 8'hA2;
                    16'hDE3D: data_out = 8'hA1;
                    16'hDE3E: data_out = 8'hA0;
                    16'hDE3F: data_out = 8'h9F;
                    16'hDE40: data_out = 8'h9E;
                    16'hDE41: data_out = 8'h9D;
                    16'hDE42: data_out = 8'h9C;
                    16'hDE43: data_out = 8'h9B;
                    16'hDE44: data_out = 8'h9A;
                    16'hDE45: data_out = 8'h99;
                    16'hDE46: data_out = 8'h98;
                    16'hDE47: data_out = 8'h97;
                    16'hDE48: data_out = 8'h96;
                    16'hDE49: data_out = 8'h95;
                    16'hDE4A: data_out = 8'h94;
                    16'hDE4B: data_out = 8'h93;
                    16'hDE4C: data_out = 8'h92;
                    16'hDE4D: data_out = 8'h91;
                    16'hDE4E: data_out = 8'h90;
                    16'hDE4F: data_out = 8'h8F;
                    16'hDE50: data_out = 8'h8E;
                    16'hDE51: data_out = 8'h8D;
                    16'hDE52: data_out = 8'h8C;
                    16'hDE53: data_out = 8'h8B;
                    16'hDE54: data_out = 8'h8A;
                    16'hDE55: data_out = 8'h89;
                    16'hDE56: data_out = 8'h88;
                    16'hDE57: data_out = 8'h87;
                    16'hDE58: data_out = 8'h86;
                    16'hDE59: data_out = 8'h85;
                    16'hDE5A: data_out = 8'h84;
                    16'hDE5B: data_out = 8'h83;
                    16'hDE5C: data_out = 8'h82;
                    16'hDE5D: data_out = 8'h81;
                    16'hDE5E: data_out = 8'h0;
                    16'hDE5F: data_out = 8'h1;
                    16'hDE60: data_out = 8'h2;
                    16'hDE61: data_out = 8'h3;
                    16'hDE62: data_out = 8'h4;
                    16'hDE63: data_out = 8'h5;
                    16'hDE64: data_out = 8'h6;
                    16'hDE65: data_out = 8'h7;
                    16'hDE66: data_out = 8'h8;
                    16'hDE67: data_out = 8'h9;
                    16'hDE68: data_out = 8'hA;
                    16'hDE69: data_out = 8'hB;
                    16'hDE6A: data_out = 8'hC;
                    16'hDE6B: data_out = 8'hD;
                    16'hDE6C: data_out = 8'hE;
                    16'hDE6D: data_out = 8'hF;
                    16'hDE6E: data_out = 8'h10;
                    16'hDE6F: data_out = 8'h11;
                    16'hDE70: data_out = 8'h12;
                    16'hDE71: data_out = 8'h13;
                    16'hDE72: data_out = 8'h14;
                    16'hDE73: data_out = 8'h15;
                    16'hDE74: data_out = 8'h16;
                    16'hDE75: data_out = 8'h17;
                    16'hDE76: data_out = 8'h18;
                    16'hDE77: data_out = 8'h19;
                    16'hDE78: data_out = 8'h1A;
                    16'hDE79: data_out = 8'h1B;
                    16'hDE7A: data_out = 8'h1C;
                    16'hDE7B: data_out = 8'h1D;
                    16'hDE7C: data_out = 8'h1E;
                    16'hDE7D: data_out = 8'h1F;
                    16'hDE7E: data_out = 8'h20;
                    16'hDE7F: data_out = 8'h21;
                    16'hDE80: data_out = 8'hDE;
                    16'hDE81: data_out = 8'hDF;
                    16'hDE82: data_out = 8'hE0;
                    16'hDE83: data_out = 8'hE1;
                    16'hDE84: data_out = 8'hE2;
                    16'hDE85: data_out = 8'hE3;
                    16'hDE86: data_out = 8'hE4;
                    16'hDE87: data_out = 8'hE5;
                    16'hDE88: data_out = 8'hE6;
                    16'hDE89: data_out = 8'hE7;
                    16'hDE8A: data_out = 8'hE8;
                    16'hDE8B: data_out = 8'hE9;
                    16'hDE8C: data_out = 8'hEA;
                    16'hDE8D: data_out = 8'hEB;
                    16'hDE8E: data_out = 8'hEC;
                    16'hDE8F: data_out = 8'hED;
                    16'hDE90: data_out = 8'hEE;
                    16'hDE91: data_out = 8'hEF;
                    16'hDE92: data_out = 8'hF0;
                    16'hDE93: data_out = 8'hF1;
                    16'hDE94: data_out = 8'hF2;
                    16'hDE95: data_out = 8'hF3;
                    16'hDE96: data_out = 8'hF4;
                    16'hDE97: data_out = 8'hF5;
                    16'hDE98: data_out = 8'hF6;
                    16'hDE99: data_out = 8'hF7;
                    16'hDE9A: data_out = 8'hF8;
                    16'hDE9B: data_out = 8'hF9;
                    16'hDE9C: data_out = 8'hFA;
                    16'hDE9D: data_out = 8'hFB;
                    16'hDE9E: data_out = 8'hFC;
                    16'hDE9F: data_out = 8'hFD;
                    16'hDEA0: data_out = 8'hFE;
                    16'hDEA1: data_out = 8'hFF;
                    16'hDEA2: data_out = 8'h80;
                    16'hDEA3: data_out = 8'h81;
                    16'hDEA4: data_out = 8'h82;
                    16'hDEA5: data_out = 8'h83;
                    16'hDEA6: data_out = 8'h84;
                    16'hDEA7: data_out = 8'h85;
                    16'hDEA8: data_out = 8'h86;
                    16'hDEA9: data_out = 8'h87;
                    16'hDEAA: data_out = 8'h88;
                    16'hDEAB: data_out = 8'h89;
                    16'hDEAC: data_out = 8'h8A;
                    16'hDEAD: data_out = 8'h8B;
                    16'hDEAE: data_out = 8'h8C;
                    16'hDEAF: data_out = 8'h8D;
                    16'hDEB0: data_out = 8'h8E;
                    16'hDEB1: data_out = 8'h8F;
                    16'hDEB2: data_out = 8'h90;
                    16'hDEB3: data_out = 8'h91;
                    16'hDEB4: data_out = 8'h92;
                    16'hDEB5: data_out = 8'h93;
                    16'hDEB6: data_out = 8'h94;
                    16'hDEB7: data_out = 8'h95;
                    16'hDEB8: data_out = 8'h96;
                    16'hDEB9: data_out = 8'h97;
                    16'hDEBA: data_out = 8'h98;
                    16'hDEBB: data_out = 8'h99;
                    16'hDEBC: data_out = 8'h9A;
                    16'hDEBD: data_out = 8'h9B;
                    16'hDEBE: data_out = 8'h9C;
                    16'hDEBF: data_out = 8'h9D;
                    16'hDEC0: data_out = 8'h9E;
                    16'hDEC1: data_out = 8'h9F;
                    16'hDEC2: data_out = 8'hA0;
                    16'hDEC3: data_out = 8'hA1;
                    16'hDEC4: data_out = 8'hA2;
                    16'hDEC5: data_out = 8'hA3;
                    16'hDEC6: data_out = 8'hA4;
                    16'hDEC7: data_out = 8'hA5;
                    16'hDEC8: data_out = 8'hA6;
                    16'hDEC9: data_out = 8'hA7;
                    16'hDECA: data_out = 8'hA8;
                    16'hDECB: data_out = 8'hA9;
                    16'hDECC: data_out = 8'hAA;
                    16'hDECD: data_out = 8'hAB;
                    16'hDECE: data_out = 8'hAC;
                    16'hDECF: data_out = 8'hAD;
                    16'hDED0: data_out = 8'hAE;
                    16'hDED1: data_out = 8'hAF;
                    16'hDED2: data_out = 8'hB0;
                    16'hDED3: data_out = 8'hB1;
                    16'hDED4: data_out = 8'hB2;
                    16'hDED5: data_out = 8'hB3;
                    16'hDED6: data_out = 8'hB4;
                    16'hDED7: data_out = 8'hB5;
                    16'hDED8: data_out = 8'hB6;
                    16'hDED9: data_out = 8'hB7;
                    16'hDEDA: data_out = 8'hB8;
                    16'hDEDB: data_out = 8'hB9;
                    16'hDEDC: data_out = 8'hBA;
                    16'hDEDD: data_out = 8'hBB;
                    16'hDEDE: data_out = 8'hBC;
                    16'hDEDF: data_out = 8'hBD;
                    16'hDEE0: data_out = 8'hBE;
                    16'hDEE1: data_out = 8'hBF;
                    16'hDEE2: data_out = 8'hC0;
                    16'hDEE3: data_out = 8'hC1;
                    16'hDEE4: data_out = 8'hC2;
                    16'hDEE5: data_out = 8'hC3;
                    16'hDEE6: data_out = 8'hC4;
                    16'hDEE7: data_out = 8'hC5;
                    16'hDEE8: data_out = 8'hC6;
                    16'hDEE9: data_out = 8'hC7;
                    16'hDEEA: data_out = 8'hC8;
                    16'hDEEB: data_out = 8'hC9;
                    16'hDEEC: data_out = 8'hCA;
                    16'hDEED: data_out = 8'hCB;
                    16'hDEEE: data_out = 8'hCC;
                    16'hDEEF: data_out = 8'hCD;
                    16'hDEF0: data_out = 8'hCE;
                    16'hDEF1: data_out = 8'hCF;
                    16'hDEF2: data_out = 8'hD0;
                    16'hDEF3: data_out = 8'hD1;
                    16'hDEF4: data_out = 8'hD2;
                    16'hDEF5: data_out = 8'hD3;
                    16'hDEF6: data_out = 8'hD4;
                    16'hDEF7: data_out = 8'hD5;
                    16'hDEF8: data_out = 8'hD6;
                    16'hDEF9: data_out = 8'hD7;
                    16'hDEFA: data_out = 8'hD8;
                    16'hDEFB: data_out = 8'hD9;
                    16'hDEFC: data_out = 8'hDA;
                    16'hDEFD: data_out = 8'hDB;
                    16'hDEFE: data_out = 8'hDC;
                    16'hDEFF: data_out = 8'hDD;
                    16'hDF00: data_out = 8'hDF;
                    16'hDF01: data_out = 8'hDE;
                    16'hDF02: data_out = 8'hDD;
                    16'hDF03: data_out = 8'hDC;
                    16'hDF04: data_out = 8'hDB;
                    16'hDF05: data_out = 8'hDA;
                    16'hDF06: data_out = 8'hD9;
                    16'hDF07: data_out = 8'hD8;
                    16'hDF08: data_out = 8'hD7;
                    16'hDF09: data_out = 8'hD6;
                    16'hDF0A: data_out = 8'hD5;
                    16'hDF0B: data_out = 8'hD4;
                    16'hDF0C: data_out = 8'hD3;
                    16'hDF0D: data_out = 8'hD2;
                    16'hDF0E: data_out = 8'hD1;
                    16'hDF0F: data_out = 8'hD0;
                    16'hDF10: data_out = 8'hCF;
                    16'hDF11: data_out = 8'hCE;
                    16'hDF12: data_out = 8'hCD;
                    16'hDF13: data_out = 8'hCC;
                    16'hDF14: data_out = 8'hCB;
                    16'hDF15: data_out = 8'hCA;
                    16'hDF16: data_out = 8'hC9;
                    16'hDF17: data_out = 8'hC8;
                    16'hDF18: data_out = 8'hC7;
                    16'hDF19: data_out = 8'hC6;
                    16'hDF1A: data_out = 8'hC5;
                    16'hDF1B: data_out = 8'hC4;
                    16'hDF1C: data_out = 8'hC3;
                    16'hDF1D: data_out = 8'hC2;
                    16'hDF1E: data_out = 8'hC1;
                    16'hDF1F: data_out = 8'hC0;
                    16'hDF20: data_out = 8'hBF;
                    16'hDF21: data_out = 8'hBE;
                    16'hDF22: data_out = 8'hBD;
                    16'hDF23: data_out = 8'hBC;
                    16'hDF24: data_out = 8'hBB;
                    16'hDF25: data_out = 8'hBA;
                    16'hDF26: data_out = 8'hB9;
                    16'hDF27: data_out = 8'hB8;
                    16'hDF28: data_out = 8'hB7;
                    16'hDF29: data_out = 8'hB6;
                    16'hDF2A: data_out = 8'hB5;
                    16'hDF2B: data_out = 8'hB4;
                    16'hDF2C: data_out = 8'hB3;
                    16'hDF2D: data_out = 8'hB2;
                    16'hDF2E: data_out = 8'hB1;
                    16'hDF2F: data_out = 8'hB0;
                    16'hDF30: data_out = 8'hAF;
                    16'hDF31: data_out = 8'hAE;
                    16'hDF32: data_out = 8'hAD;
                    16'hDF33: data_out = 8'hAC;
                    16'hDF34: data_out = 8'hAB;
                    16'hDF35: data_out = 8'hAA;
                    16'hDF36: data_out = 8'hA9;
                    16'hDF37: data_out = 8'hA8;
                    16'hDF38: data_out = 8'hA7;
                    16'hDF39: data_out = 8'hA6;
                    16'hDF3A: data_out = 8'hA5;
                    16'hDF3B: data_out = 8'hA4;
                    16'hDF3C: data_out = 8'hA3;
                    16'hDF3D: data_out = 8'hA2;
                    16'hDF3E: data_out = 8'hA1;
                    16'hDF3F: data_out = 8'hA0;
                    16'hDF40: data_out = 8'h9F;
                    16'hDF41: data_out = 8'h9E;
                    16'hDF42: data_out = 8'h9D;
                    16'hDF43: data_out = 8'h9C;
                    16'hDF44: data_out = 8'h9B;
                    16'hDF45: data_out = 8'h9A;
                    16'hDF46: data_out = 8'h99;
                    16'hDF47: data_out = 8'h98;
                    16'hDF48: data_out = 8'h97;
                    16'hDF49: data_out = 8'h96;
                    16'hDF4A: data_out = 8'h95;
                    16'hDF4B: data_out = 8'h94;
                    16'hDF4C: data_out = 8'h93;
                    16'hDF4D: data_out = 8'h92;
                    16'hDF4E: data_out = 8'h91;
                    16'hDF4F: data_out = 8'h90;
                    16'hDF50: data_out = 8'h8F;
                    16'hDF51: data_out = 8'h8E;
                    16'hDF52: data_out = 8'h8D;
                    16'hDF53: data_out = 8'h8C;
                    16'hDF54: data_out = 8'h8B;
                    16'hDF55: data_out = 8'h8A;
                    16'hDF56: data_out = 8'h89;
                    16'hDF57: data_out = 8'h88;
                    16'hDF58: data_out = 8'h87;
                    16'hDF59: data_out = 8'h86;
                    16'hDF5A: data_out = 8'h85;
                    16'hDF5B: data_out = 8'h84;
                    16'hDF5C: data_out = 8'h83;
                    16'hDF5D: data_out = 8'h82;
                    16'hDF5E: data_out = 8'h81;
                    16'hDF5F: data_out = 8'h0;
                    16'hDF60: data_out = 8'h1;
                    16'hDF61: data_out = 8'h2;
                    16'hDF62: data_out = 8'h3;
                    16'hDF63: data_out = 8'h4;
                    16'hDF64: data_out = 8'h5;
                    16'hDF65: data_out = 8'h6;
                    16'hDF66: data_out = 8'h7;
                    16'hDF67: data_out = 8'h8;
                    16'hDF68: data_out = 8'h9;
                    16'hDF69: data_out = 8'hA;
                    16'hDF6A: data_out = 8'hB;
                    16'hDF6B: data_out = 8'hC;
                    16'hDF6C: data_out = 8'hD;
                    16'hDF6D: data_out = 8'hE;
                    16'hDF6E: data_out = 8'hF;
                    16'hDF6F: data_out = 8'h10;
                    16'hDF70: data_out = 8'h11;
                    16'hDF71: data_out = 8'h12;
                    16'hDF72: data_out = 8'h13;
                    16'hDF73: data_out = 8'h14;
                    16'hDF74: data_out = 8'h15;
                    16'hDF75: data_out = 8'h16;
                    16'hDF76: data_out = 8'h17;
                    16'hDF77: data_out = 8'h18;
                    16'hDF78: data_out = 8'h19;
                    16'hDF79: data_out = 8'h1A;
                    16'hDF7A: data_out = 8'h1B;
                    16'hDF7B: data_out = 8'h1C;
                    16'hDF7C: data_out = 8'h1D;
                    16'hDF7D: data_out = 8'h1E;
                    16'hDF7E: data_out = 8'h1F;
                    16'hDF7F: data_out = 8'h20;
                    16'hDF80: data_out = 8'hDF;
                    16'hDF81: data_out = 8'hE0;
                    16'hDF82: data_out = 8'hE1;
                    16'hDF83: data_out = 8'hE2;
                    16'hDF84: data_out = 8'hE3;
                    16'hDF85: data_out = 8'hE4;
                    16'hDF86: data_out = 8'hE5;
                    16'hDF87: data_out = 8'hE6;
                    16'hDF88: data_out = 8'hE7;
                    16'hDF89: data_out = 8'hE8;
                    16'hDF8A: data_out = 8'hE9;
                    16'hDF8B: data_out = 8'hEA;
                    16'hDF8C: data_out = 8'hEB;
                    16'hDF8D: data_out = 8'hEC;
                    16'hDF8E: data_out = 8'hED;
                    16'hDF8F: data_out = 8'hEE;
                    16'hDF90: data_out = 8'hEF;
                    16'hDF91: data_out = 8'hF0;
                    16'hDF92: data_out = 8'hF1;
                    16'hDF93: data_out = 8'hF2;
                    16'hDF94: data_out = 8'hF3;
                    16'hDF95: data_out = 8'hF4;
                    16'hDF96: data_out = 8'hF5;
                    16'hDF97: data_out = 8'hF6;
                    16'hDF98: data_out = 8'hF7;
                    16'hDF99: data_out = 8'hF8;
                    16'hDF9A: data_out = 8'hF9;
                    16'hDF9B: data_out = 8'hFA;
                    16'hDF9C: data_out = 8'hFB;
                    16'hDF9D: data_out = 8'hFC;
                    16'hDF9E: data_out = 8'hFD;
                    16'hDF9F: data_out = 8'hFE;
                    16'hDFA0: data_out = 8'hFF;
                    16'hDFA1: data_out = 8'h80;
                    16'hDFA2: data_out = 8'h81;
                    16'hDFA3: data_out = 8'h82;
                    16'hDFA4: data_out = 8'h83;
                    16'hDFA5: data_out = 8'h84;
                    16'hDFA6: data_out = 8'h85;
                    16'hDFA7: data_out = 8'h86;
                    16'hDFA8: data_out = 8'h87;
                    16'hDFA9: data_out = 8'h88;
                    16'hDFAA: data_out = 8'h89;
                    16'hDFAB: data_out = 8'h8A;
                    16'hDFAC: data_out = 8'h8B;
                    16'hDFAD: data_out = 8'h8C;
                    16'hDFAE: data_out = 8'h8D;
                    16'hDFAF: data_out = 8'h8E;
                    16'hDFB0: data_out = 8'h8F;
                    16'hDFB1: data_out = 8'h90;
                    16'hDFB2: data_out = 8'h91;
                    16'hDFB3: data_out = 8'h92;
                    16'hDFB4: data_out = 8'h93;
                    16'hDFB5: data_out = 8'h94;
                    16'hDFB6: data_out = 8'h95;
                    16'hDFB7: data_out = 8'h96;
                    16'hDFB8: data_out = 8'h97;
                    16'hDFB9: data_out = 8'h98;
                    16'hDFBA: data_out = 8'h99;
                    16'hDFBB: data_out = 8'h9A;
                    16'hDFBC: data_out = 8'h9B;
                    16'hDFBD: data_out = 8'h9C;
                    16'hDFBE: data_out = 8'h9D;
                    16'hDFBF: data_out = 8'h9E;
                    16'hDFC0: data_out = 8'h9F;
                    16'hDFC1: data_out = 8'hA0;
                    16'hDFC2: data_out = 8'hA1;
                    16'hDFC3: data_out = 8'hA2;
                    16'hDFC4: data_out = 8'hA3;
                    16'hDFC5: data_out = 8'hA4;
                    16'hDFC6: data_out = 8'hA5;
                    16'hDFC7: data_out = 8'hA6;
                    16'hDFC8: data_out = 8'hA7;
                    16'hDFC9: data_out = 8'hA8;
                    16'hDFCA: data_out = 8'hA9;
                    16'hDFCB: data_out = 8'hAA;
                    16'hDFCC: data_out = 8'hAB;
                    16'hDFCD: data_out = 8'hAC;
                    16'hDFCE: data_out = 8'hAD;
                    16'hDFCF: data_out = 8'hAE;
                    16'hDFD0: data_out = 8'hAF;
                    16'hDFD1: data_out = 8'hB0;
                    16'hDFD2: data_out = 8'hB1;
                    16'hDFD3: data_out = 8'hB2;
                    16'hDFD4: data_out = 8'hB3;
                    16'hDFD5: data_out = 8'hB4;
                    16'hDFD6: data_out = 8'hB5;
                    16'hDFD7: data_out = 8'hB6;
                    16'hDFD8: data_out = 8'hB7;
                    16'hDFD9: data_out = 8'hB8;
                    16'hDFDA: data_out = 8'hB9;
                    16'hDFDB: data_out = 8'hBA;
                    16'hDFDC: data_out = 8'hBB;
                    16'hDFDD: data_out = 8'hBC;
                    16'hDFDE: data_out = 8'hBD;
                    16'hDFDF: data_out = 8'hBE;
                    16'hDFE0: data_out = 8'hBF;
                    16'hDFE1: data_out = 8'hC0;
                    16'hDFE2: data_out = 8'hC1;
                    16'hDFE3: data_out = 8'hC2;
                    16'hDFE4: data_out = 8'hC3;
                    16'hDFE5: data_out = 8'hC4;
                    16'hDFE6: data_out = 8'hC5;
                    16'hDFE7: data_out = 8'hC6;
                    16'hDFE8: data_out = 8'hC7;
                    16'hDFE9: data_out = 8'hC8;
                    16'hDFEA: data_out = 8'hC9;
                    16'hDFEB: data_out = 8'hCA;
                    16'hDFEC: data_out = 8'hCB;
                    16'hDFED: data_out = 8'hCC;
                    16'hDFEE: data_out = 8'hCD;
                    16'hDFEF: data_out = 8'hCE;
                    16'hDFF0: data_out = 8'hCF;
                    16'hDFF1: data_out = 8'hD0;
                    16'hDFF2: data_out = 8'hD1;
                    16'hDFF3: data_out = 8'hD2;
                    16'hDFF4: data_out = 8'hD3;
                    16'hDFF5: data_out = 8'hD4;
                    16'hDFF6: data_out = 8'hD5;
                    16'hDFF7: data_out = 8'hD6;
                    16'hDFF8: data_out = 8'hD7;
                    16'hDFF9: data_out = 8'hD8;
                    16'hDFFA: data_out = 8'hD9;
                    16'hDFFB: data_out = 8'hDA;
                    16'hDFFC: data_out = 8'hDB;
                    16'hDFFD: data_out = 8'hDC;
                    16'hDFFE: data_out = 8'hDD;
                    16'hDFFF: data_out = 8'hDE;
                    16'hE000: data_out = 8'hE0;
                    16'hE001: data_out = 8'hDF;
                    16'hE002: data_out = 8'hDE;
                    16'hE003: data_out = 8'hDD;
                    16'hE004: data_out = 8'hDC;
                    16'hE005: data_out = 8'hDB;
                    16'hE006: data_out = 8'hDA;
                    16'hE007: data_out = 8'hD9;
                    16'hE008: data_out = 8'hD8;
                    16'hE009: data_out = 8'hD7;
                    16'hE00A: data_out = 8'hD6;
                    16'hE00B: data_out = 8'hD5;
                    16'hE00C: data_out = 8'hD4;
                    16'hE00D: data_out = 8'hD3;
                    16'hE00E: data_out = 8'hD2;
                    16'hE00F: data_out = 8'hD1;
                    16'hE010: data_out = 8'hD0;
                    16'hE011: data_out = 8'hCF;
                    16'hE012: data_out = 8'hCE;
                    16'hE013: data_out = 8'hCD;
                    16'hE014: data_out = 8'hCC;
                    16'hE015: data_out = 8'hCB;
                    16'hE016: data_out = 8'hCA;
                    16'hE017: data_out = 8'hC9;
                    16'hE018: data_out = 8'hC8;
                    16'hE019: data_out = 8'hC7;
                    16'hE01A: data_out = 8'hC6;
                    16'hE01B: data_out = 8'hC5;
                    16'hE01C: data_out = 8'hC4;
                    16'hE01D: data_out = 8'hC3;
                    16'hE01E: data_out = 8'hC2;
                    16'hE01F: data_out = 8'hC1;
                    16'hE020: data_out = 8'hC0;
                    16'hE021: data_out = 8'hBF;
                    16'hE022: data_out = 8'hBE;
                    16'hE023: data_out = 8'hBD;
                    16'hE024: data_out = 8'hBC;
                    16'hE025: data_out = 8'hBB;
                    16'hE026: data_out = 8'hBA;
                    16'hE027: data_out = 8'hB9;
                    16'hE028: data_out = 8'hB8;
                    16'hE029: data_out = 8'hB7;
                    16'hE02A: data_out = 8'hB6;
                    16'hE02B: data_out = 8'hB5;
                    16'hE02C: data_out = 8'hB4;
                    16'hE02D: data_out = 8'hB3;
                    16'hE02E: data_out = 8'hB2;
                    16'hE02F: data_out = 8'hB1;
                    16'hE030: data_out = 8'hB0;
                    16'hE031: data_out = 8'hAF;
                    16'hE032: data_out = 8'hAE;
                    16'hE033: data_out = 8'hAD;
                    16'hE034: data_out = 8'hAC;
                    16'hE035: data_out = 8'hAB;
                    16'hE036: data_out = 8'hAA;
                    16'hE037: data_out = 8'hA9;
                    16'hE038: data_out = 8'hA8;
                    16'hE039: data_out = 8'hA7;
                    16'hE03A: data_out = 8'hA6;
                    16'hE03B: data_out = 8'hA5;
                    16'hE03C: data_out = 8'hA4;
                    16'hE03D: data_out = 8'hA3;
                    16'hE03E: data_out = 8'hA2;
                    16'hE03F: data_out = 8'hA1;
                    16'hE040: data_out = 8'hA0;
                    16'hE041: data_out = 8'h9F;
                    16'hE042: data_out = 8'h9E;
                    16'hE043: data_out = 8'h9D;
                    16'hE044: data_out = 8'h9C;
                    16'hE045: data_out = 8'h9B;
                    16'hE046: data_out = 8'h9A;
                    16'hE047: data_out = 8'h99;
                    16'hE048: data_out = 8'h98;
                    16'hE049: data_out = 8'h97;
                    16'hE04A: data_out = 8'h96;
                    16'hE04B: data_out = 8'h95;
                    16'hE04C: data_out = 8'h94;
                    16'hE04D: data_out = 8'h93;
                    16'hE04E: data_out = 8'h92;
                    16'hE04F: data_out = 8'h91;
                    16'hE050: data_out = 8'h90;
                    16'hE051: data_out = 8'h8F;
                    16'hE052: data_out = 8'h8E;
                    16'hE053: data_out = 8'h8D;
                    16'hE054: data_out = 8'h8C;
                    16'hE055: data_out = 8'h8B;
                    16'hE056: data_out = 8'h8A;
                    16'hE057: data_out = 8'h89;
                    16'hE058: data_out = 8'h88;
                    16'hE059: data_out = 8'h87;
                    16'hE05A: data_out = 8'h86;
                    16'hE05B: data_out = 8'h85;
                    16'hE05C: data_out = 8'h84;
                    16'hE05D: data_out = 8'h83;
                    16'hE05E: data_out = 8'h82;
                    16'hE05F: data_out = 8'h81;
                    16'hE060: data_out = 8'h0;
                    16'hE061: data_out = 8'h1;
                    16'hE062: data_out = 8'h2;
                    16'hE063: data_out = 8'h3;
                    16'hE064: data_out = 8'h4;
                    16'hE065: data_out = 8'h5;
                    16'hE066: data_out = 8'h6;
                    16'hE067: data_out = 8'h7;
                    16'hE068: data_out = 8'h8;
                    16'hE069: data_out = 8'h9;
                    16'hE06A: data_out = 8'hA;
                    16'hE06B: data_out = 8'hB;
                    16'hE06C: data_out = 8'hC;
                    16'hE06D: data_out = 8'hD;
                    16'hE06E: data_out = 8'hE;
                    16'hE06F: data_out = 8'hF;
                    16'hE070: data_out = 8'h10;
                    16'hE071: data_out = 8'h11;
                    16'hE072: data_out = 8'h12;
                    16'hE073: data_out = 8'h13;
                    16'hE074: data_out = 8'h14;
                    16'hE075: data_out = 8'h15;
                    16'hE076: data_out = 8'h16;
                    16'hE077: data_out = 8'h17;
                    16'hE078: data_out = 8'h18;
                    16'hE079: data_out = 8'h19;
                    16'hE07A: data_out = 8'h1A;
                    16'hE07B: data_out = 8'h1B;
                    16'hE07C: data_out = 8'h1C;
                    16'hE07D: data_out = 8'h1D;
                    16'hE07E: data_out = 8'h1E;
                    16'hE07F: data_out = 8'h1F;
                    16'hE080: data_out = 8'hE0;
                    16'hE081: data_out = 8'hE1;
                    16'hE082: data_out = 8'hE2;
                    16'hE083: data_out = 8'hE3;
                    16'hE084: data_out = 8'hE4;
                    16'hE085: data_out = 8'hE5;
                    16'hE086: data_out = 8'hE6;
                    16'hE087: data_out = 8'hE7;
                    16'hE088: data_out = 8'hE8;
                    16'hE089: data_out = 8'hE9;
                    16'hE08A: data_out = 8'hEA;
                    16'hE08B: data_out = 8'hEB;
                    16'hE08C: data_out = 8'hEC;
                    16'hE08D: data_out = 8'hED;
                    16'hE08E: data_out = 8'hEE;
                    16'hE08F: data_out = 8'hEF;
                    16'hE090: data_out = 8'hF0;
                    16'hE091: data_out = 8'hF1;
                    16'hE092: data_out = 8'hF2;
                    16'hE093: data_out = 8'hF3;
                    16'hE094: data_out = 8'hF4;
                    16'hE095: data_out = 8'hF5;
                    16'hE096: data_out = 8'hF6;
                    16'hE097: data_out = 8'hF7;
                    16'hE098: data_out = 8'hF8;
                    16'hE099: data_out = 8'hF9;
                    16'hE09A: data_out = 8'hFA;
                    16'hE09B: data_out = 8'hFB;
                    16'hE09C: data_out = 8'hFC;
                    16'hE09D: data_out = 8'hFD;
                    16'hE09E: data_out = 8'hFE;
                    16'hE09F: data_out = 8'hFF;
                    16'hE0A0: data_out = 8'h80;
                    16'hE0A1: data_out = 8'h81;
                    16'hE0A2: data_out = 8'h82;
                    16'hE0A3: data_out = 8'h83;
                    16'hE0A4: data_out = 8'h84;
                    16'hE0A5: data_out = 8'h85;
                    16'hE0A6: data_out = 8'h86;
                    16'hE0A7: data_out = 8'h87;
                    16'hE0A8: data_out = 8'h88;
                    16'hE0A9: data_out = 8'h89;
                    16'hE0AA: data_out = 8'h8A;
                    16'hE0AB: data_out = 8'h8B;
                    16'hE0AC: data_out = 8'h8C;
                    16'hE0AD: data_out = 8'h8D;
                    16'hE0AE: data_out = 8'h8E;
                    16'hE0AF: data_out = 8'h8F;
                    16'hE0B0: data_out = 8'h90;
                    16'hE0B1: data_out = 8'h91;
                    16'hE0B2: data_out = 8'h92;
                    16'hE0B3: data_out = 8'h93;
                    16'hE0B4: data_out = 8'h94;
                    16'hE0B5: data_out = 8'h95;
                    16'hE0B6: data_out = 8'h96;
                    16'hE0B7: data_out = 8'h97;
                    16'hE0B8: data_out = 8'h98;
                    16'hE0B9: data_out = 8'h99;
                    16'hE0BA: data_out = 8'h9A;
                    16'hE0BB: data_out = 8'h9B;
                    16'hE0BC: data_out = 8'h9C;
                    16'hE0BD: data_out = 8'h9D;
                    16'hE0BE: data_out = 8'h9E;
                    16'hE0BF: data_out = 8'h9F;
                    16'hE0C0: data_out = 8'hA0;
                    16'hE0C1: data_out = 8'hA1;
                    16'hE0C2: data_out = 8'hA2;
                    16'hE0C3: data_out = 8'hA3;
                    16'hE0C4: data_out = 8'hA4;
                    16'hE0C5: data_out = 8'hA5;
                    16'hE0C6: data_out = 8'hA6;
                    16'hE0C7: data_out = 8'hA7;
                    16'hE0C8: data_out = 8'hA8;
                    16'hE0C9: data_out = 8'hA9;
                    16'hE0CA: data_out = 8'hAA;
                    16'hE0CB: data_out = 8'hAB;
                    16'hE0CC: data_out = 8'hAC;
                    16'hE0CD: data_out = 8'hAD;
                    16'hE0CE: data_out = 8'hAE;
                    16'hE0CF: data_out = 8'hAF;
                    16'hE0D0: data_out = 8'hB0;
                    16'hE0D1: data_out = 8'hB1;
                    16'hE0D2: data_out = 8'hB2;
                    16'hE0D3: data_out = 8'hB3;
                    16'hE0D4: data_out = 8'hB4;
                    16'hE0D5: data_out = 8'hB5;
                    16'hE0D6: data_out = 8'hB6;
                    16'hE0D7: data_out = 8'hB7;
                    16'hE0D8: data_out = 8'hB8;
                    16'hE0D9: data_out = 8'hB9;
                    16'hE0DA: data_out = 8'hBA;
                    16'hE0DB: data_out = 8'hBB;
                    16'hE0DC: data_out = 8'hBC;
                    16'hE0DD: data_out = 8'hBD;
                    16'hE0DE: data_out = 8'hBE;
                    16'hE0DF: data_out = 8'hBF;
                    16'hE0E0: data_out = 8'hC0;
                    16'hE0E1: data_out = 8'hC1;
                    16'hE0E2: data_out = 8'hC2;
                    16'hE0E3: data_out = 8'hC3;
                    16'hE0E4: data_out = 8'hC4;
                    16'hE0E5: data_out = 8'hC5;
                    16'hE0E6: data_out = 8'hC6;
                    16'hE0E7: data_out = 8'hC7;
                    16'hE0E8: data_out = 8'hC8;
                    16'hE0E9: data_out = 8'hC9;
                    16'hE0EA: data_out = 8'hCA;
                    16'hE0EB: data_out = 8'hCB;
                    16'hE0EC: data_out = 8'hCC;
                    16'hE0ED: data_out = 8'hCD;
                    16'hE0EE: data_out = 8'hCE;
                    16'hE0EF: data_out = 8'hCF;
                    16'hE0F0: data_out = 8'hD0;
                    16'hE0F1: data_out = 8'hD1;
                    16'hE0F2: data_out = 8'hD2;
                    16'hE0F3: data_out = 8'hD3;
                    16'hE0F4: data_out = 8'hD4;
                    16'hE0F5: data_out = 8'hD5;
                    16'hE0F6: data_out = 8'hD6;
                    16'hE0F7: data_out = 8'hD7;
                    16'hE0F8: data_out = 8'hD8;
                    16'hE0F9: data_out = 8'hD9;
                    16'hE0FA: data_out = 8'hDA;
                    16'hE0FB: data_out = 8'hDB;
                    16'hE0FC: data_out = 8'hDC;
                    16'hE0FD: data_out = 8'hDD;
                    16'hE0FE: data_out = 8'hDE;
                    16'hE0FF: data_out = 8'hDF;
                    16'hE100: data_out = 8'hE1;
                    16'hE101: data_out = 8'hE0;
                    16'hE102: data_out = 8'hDF;
                    16'hE103: data_out = 8'hDE;
                    16'hE104: data_out = 8'hDD;
                    16'hE105: data_out = 8'hDC;
                    16'hE106: data_out = 8'hDB;
                    16'hE107: data_out = 8'hDA;
                    16'hE108: data_out = 8'hD9;
                    16'hE109: data_out = 8'hD8;
                    16'hE10A: data_out = 8'hD7;
                    16'hE10B: data_out = 8'hD6;
                    16'hE10C: data_out = 8'hD5;
                    16'hE10D: data_out = 8'hD4;
                    16'hE10E: data_out = 8'hD3;
                    16'hE10F: data_out = 8'hD2;
                    16'hE110: data_out = 8'hD1;
                    16'hE111: data_out = 8'hD0;
                    16'hE112: data_out = 8'hCF;
                    16'hE113: data_out = 8'hCE;
                    16'hE114: data_out = 8'hCD;
                    16'hE115: data_out = 8'hCC;
                    16'hE116: data_out = 8'hCB;
                    16'hE117: data_out = 8'hCA;
                    16'hE118: data_out = 8'hC9;
                    16'hE119: data_out = 8'hC8;
                    16'hE11A: data_out = 8'hC7;
                    16'hE11B: data_out = 8'hC6;
                    16'hE11C: data_out = 8'hC5;
                    16'hE11D: data_out = 8'hC4;
                    16'hE11E: data_out = 8'hC3;
                    16'hE11F: data_out = 8'hC2;
                    16'hE120: data_out = 8'hC1;
                    16'hE121: data_out = 8'hC0;
                    16'hE122: data_out = 8'hBF;
                    16'hE123: data_out = 8'hBE;
                    16'hE124: data_out = 8'hBD;
                    16'hE125: data_out = 8'hBC;
                    16'hE126: data_out = 8'hBB;
                    16'hE127: data_out = 8'hBA;
                    16'hE128: data_out = 8'hB9;
                    16'hE129: data_out = 8'hB8;
                    16'hE12A: data_out = 8'hB7;
                    16'hE12B: data_out = 8'hB6;
                    16'hE12C: data_out = 8'hB5;
                    16'hE12D: data_out = 8'hB4;
                    16'hE12E: data_out = 8'hB3;
                    16'hE12F: data_out = 8'hB2;
                    16'hE130: data_out = 8'hB1;
                    16'hE131: data_out = 8'hB0;
                    16'hE132: data_out = 8'hAF;
                    16'hE133: data_out = 8'hAE;
                    16'hE134: data_out = 8'hAD;
                    16'hE135: data_out = 8'hAC;
                    16'hE136: data_out = 8'hAB;
                    16'hE137: data_out = 8'hAA;
                    16'hE138: data_out = 8'hA9;
                    16'hE139: data_out = 8'hA8;
                    16'hE13A: data_out = 8'hA7;
                    16'hE13B: data_out = 8'hA6;
                    16'hE13C: data_out = 8'hA5;
                    16'hE13D: data_out = 8'hA4;
                    16'hE13E: data_out = 8'hA3;
                    16'hE13F: data_out = 8'hA2;
                    16'hE140: data_out = 8'hA1;
                    16'hE141: data_out = 8'hA0;
                    16'hE142: data_out = 8'h9F;
                    16'hE143: data_out = 8'h9E;
                    16'hE144: data_out = 8'h9D;
                    16'hE145: data_out = 8'h9C;
                    16'hE146: data_out = 8'h9B;
                    16'hE147: data_out = 8'h9A;
                    16'hE148: data_out = 8'h99;
                    16'hE149: data_out = 8'h98;
                    16'hE14A: data_out = 8'h97;
                    16'hE14B: data_out = 8'h96;
                    16'hE14C: data_out = 8'h95;
                    16'hE14D: data_out = 8'h94;
                    16'hE14E: data_out = 8'h93;
                    16'hE14F: data_out = 8'h92;
                    16'hE150: data_out = 8'h91;
                    16'hE151: data_out = 8'h90;
                    16'hE152: data_out = 8'h8F;
                    16'hE153: data_out = 8'h8E;
                    16'hE154: data_out = 8'h8D;
                    16'hE155: data_out = 8'h8C;
                    16'hE156: data_out = 8'h8B;
                    16'hE157: data_out = 8'h8A;
                    16'hE158: data_out = 8'h89;
                    16'hE159: data_out = 8'h88;
                    16'hE15A: data_out = 8'h87;
                    16'hE15B: data_out = 8'h86;
                    16'hE15C: data_out = 8'h85;
                    16'hE15D: data_out = 8'h84;
                    16'hE15E: data_out = 8'h83;
                    16'hE15F: data_out = 8'h82;
                    16'hE160: data_out = 8'h81;
                    16'hE161: data_out = 8'h0;
                    16'hE162: data_out = 8'h1;
                    16'hE163: data_out = 8'h2;
                    16'hE164: data_out = 8'h3;
                    16'hE165: data_out = 8'h4;
                    16'hE166: data_out = 8'h5;
                    16'hE167: data_out = 8'h6;
                    16'hE168: data_out = 8'h7;
                    16'hE169: data_out = 8'h8;
                    16'hE16A: data_out = 8'h9;
                    16'hE16B: data_out = 8'hA;
                    16'hE16C: data_out = 8'hB;
                    16'hE16D: data_out = 8'hC;
                    16'hE16E: data_out = 8'hD;
                    16'hE16F: data_out = 8'hE;
                    16'hE170: data_out = 8'hF;
                    16'hE171: data_out = 8'h10;
                    16'hE172: data_out = 8'h11;
                    16'hE173: data_out = 8'h12;
                    16'hE174: data_out = 8'h13;
                    16'hE175: data_out = 8'h14;
                    16'hE176: data_out = 8'h15;
                    16'hE177: data_out = 8'h16;
                    16'hE178: data_out = 8'h17;
                    16'hE179: data_out = 8'h18;
                    16'hE17A: data_out = 8'h19;
                    16'hE17B: data_out = 8'h1A;
                    16'hE17C: data_out = 8'h1B;
                    16'hE17D: data_out = 8'h1C;
                    16'hE17E: data_out = 8'h1D;
                    16'hE17F: data_out = 8'h1E;
                    16'hE180: data_out = 8'hE1;
                    16'hE181: data_out = 8'hE2;
                    16'hE182: data_out = 8'hE3;
                    16'hE183: data_out = 8'hE4;
                    16'hE184: data_out = 8'hE5;
                    16'hE185: data_out = 8'hE6;
                    16'hE186: data_out = 8'hE7;
                    16'hE187: data_out = 8'hE8;
                    16'hE188: data_out = 8'hE9;
                    16'hE189: data_out = 8'hEA;
                    16'hE18A: data_out = 8'hEB;
                    16'hE18B: data_out = 8'hEC;
                    16'hE18C: data_out = 8'hED;
                    16'hE18D: data_out = 8'hEE;
                    16'hE18E: data_out = 8'hEF;
                    16'hE18F: data_out = 8'hF0;
                    16'hE190: data_out = 8'hF1;
                    16'hE191: data_out = 8'hF2;
                    16'hE192: data_out = 8'hF3;
                    16'hE193: data_out = 8'hF4;
                    16'hE194: data_out = 8'hF5;
                    16'hE195: data_out = 8'hF6;
                    16'hE196: data_out = 8'hF7;
                    16'hE197: data_out = 8'hF8;
                    16'hE198: data_out = 8'hF9;
                    16'hE199: data_out = 8'hFA;
                    16'hE19A: data_out = 8'hFB;
                    16'hE19B: data_out = 8'hFC;
                    16'hE19C: data_out = 8'hFD;
                    16'hE19D: data_out = 8'hFE;
                    16'hE19E: data_out = 8'hFF;
                    16'hE19F: data_out = 8'h80;
                    16'hE1A0: data_out = 8'h81;
                    16'hE1A1: data_out = 8'h82;
                    16'hE1A2: data_out = 8'h83;
                    16'hE1A3: data_out = 8'h84;
                    16'hE1A4: data_out = 8'h85;
                    16'hE1A5: data_out = 8'h86;
                    16'hE1A6: data_out = 8'h87;
                    16'hE1A7: data_out = 8'h88;
                    16'hE1A8: data_out = 8'h89;
                    16'hE1A9: data_out = 8'h8A;
                    16'hE1AA: data_out = 8'h8B;
                    16'hE1AB: data_out = 8'h8C;
                    16'hE1AC: data_out = 8'h8D;
                    16'hE1AD: data_out = 8'h8E;
                    16'hE1AE: data_out = 8'h8F;
                    16'hE1AF: data_out = 8'h90;
                    16'hE1B0: data_out = 8'h91;
                    16'hE1B1: data_out = 8'h92;
                    16'hE1B2: data_out = 8'h93;
                    16'hE1B3: data_out = 8'h94;
                    16'hE1B4: data_out = 8'h95;
                    16'hE1B5: data_out = 8'h96;
                    16'hE1B6: data_out = 8'h97;
                    16'hE1B7: data_out = 8'h98;
                    16'hE1B8: data_out = 8'h99;
                    16'hE1B9: data_out = 8'h9A;
                    16'hE1BA: data_out = 8'h9B;
                    16'hE1BB: data_out = 8'h9C;
                    16'hE1BC: data_out = 8'h9D;
                    16'hE1BD: data_out = 8'h9E;
                    16'hE1BE: data_out = 8'h9F;
                    16'hE1BF: data_out = 8'hA0;
                    16'hE1C0: data_out = 8'hA1;
                    16'hE1C1: data_out = 8'hA2;
                    16'hE1C2: data_out = 8'hA3;
                    16'hE1C3: data_out = 8'hA4;
                    16'hE1C4: data_out = 8'hA5;
                    16'hE1C5: data_out = 8'hA6;
                    16'hE1C6: data_out = 8'hA7;
                    16'hE1C7: data_out = 8'hA8;
                    16'hE1C8: data_out = 8'hA9;
                    16'hE1C9: data_out = 8'hAA;
                    16'hE1CA: data_out = 8'hAB;
                    16'hE1CB: data_out = 8'hAC;
                    16'hE1CC: data_out = 8'hAD;
                    16'hE1CD: data_out = 8'hAE;
                    16'hE1CE: data_out = 8'hAF;
                    16'hE1CF: data_out = 8'hB0;
                    16'hE1D0: data_out = 8'hB1;
                    16'hE1D1: data_out = 8'hB2;
                    16'hE1D2: data_out = 8'hB3;
                    16'hE1D3: data_out = 8'hB4;
                    16'hE1D4: data_out = 8'hB5;
                    16'hE1D5: data_out = 8'hB6;
                    16'hE1D6: data_out = 8'hB7;
                    16'hE1D7: data_out = 8'hB8;
                    16'hE1D8: data_out = 8'hB9;
                    16'hE1D9: data_out = 8'hBA;
                    16'hE1DA: data_out = 8'hBB;
                    16'hE1DB: data_out = 8'hBC;
                    16'hE1DC: data_out = 8'hBD;
                    16'hE1DD: data_out = 8'hBE;
                    16'hE1DE: data_out = 8'hBF;
                    16'hE1DF: data_out = 8'hC0;
                    16'hE1E0: data_out = 8'hC1;
                    16'hE1E1: data_out = 8'hC2;
                    16'hE1E2: data_out = 8'hC3;
                    16'hE1E3: data_out = 8'hC4;
                    16'hE1E4: data_out = 8'hC5;
                    16'hE1E5: data_out = 8'hC6;
                    16'hE1E6: data_out = 8'hC7;
                    16'hE1E7: data_out = 8'hC8;
                    16'hE1E8: data_out = 8'hC9;
                    16'hE1E9: data_out = 8'hCA;
                    16'hE1EA: data_out = 8'hCB;
                    16'hE1EB: data_out = 8'hCC;
                    16'hE1EC: data_out = 8'hCD;
                    16'hE1ED: data_out = 8'hCE;
                    16'hE1EE: data_out = 8'hCF;
                    16'hE1EF: data_out = 8'hD0;
                    16'hE1F0: data_out = 8'hD1;
                    16'hE1F1: data_out = 8'hD2;
                    16'hE1F2: data_out = 8'hD3;
                    16'hE1F3: data_out = 8'hD4;
                    16'hE1F4: data_out = 8'hD5;
                    16'hE1F5: data_out = 8'hD6;
                    16'hE1F6: data_out = 8'hD7;
                    16'hE1F7: data_out = 8'hD8;
                    16'hE1F8: data_out = 8'hD9;
                    16'hE1F9: data_out = 8'hDA;
                    16'hE1FA: data_out = 8'hDB;
                    16'hE1FB: data_out = 8'hDC;
                    16'hE1FC: data_out = 8'hDD;
                    16'hE1FD: data_out = 8'hDE;
                    16'hE1FE: data_out = 8'hDF;
                    16'hE1FF: data_out = 8'hE0;
                    16'hE200: data_out = 8'hE2;
                    16'hE201: data_out = 8'hE1;
                    16'hE202: data_out = 8'hE0;
                    16'hE203: data_out = 8'hDF;
                    16'hE204: data_out = 8'hDE;
                    16'hE205: data_out = 8'hDD;
                    16'hE206: data_out = 8'hDC;
                    16'hE207: data_out = 8'hDB;
                    16'hE208: data_out = 8'hDA;
                    16'hE209: data_out = 8'hD9;
                    16'hE20A: data_out = 8'hD8;
                    16'hE20B: data_out = 8'hD7;
                    16'hE20C: data_out = 8'hD6;
                    16'hE20D: data_out = 8'hD5;
                    16'hE20E: data_out = 8'hD4;
                    16'hE20F: data_out = 8'hD3;
                    16'hE210: data_out = 8'hD2;
                    16'hE211: data_out = 8'hD1;
                    16'hE212: data_out = 8'hD0;
                    16'hE213: data_out = 8'hCF;
                    16'hE214: data_out = 8'hCE;
                    16'hE215: data_out = 8'hCD;
                    16'hE216: data_out = 8'hCC;
                    16'hE217: data_out = 8'hCB;
                    16'hE218: data_out = 8'hCA;
                    16'hE219: data_out = 8'hC9;
                    16'hE21A: data_out = 8'hC8;
                    16'hE21B: data_out = 8'hC7;
                    16'hE21C: data_out = 8'hC6;
                    16'hE21D: data_out = 8'hC5;
                    16'hE21E: data_out = 8'hC4;
                    16'hE21F: data_out = 8'hC3;
                    16'hE220: data_out = 8'hC2;
                    16'hE221: data_out = 8'hC1;
                    16'hE222: data_out = 8'hC0;
                    16'hE223: data_out = 8'hBF;
                    16'hE224: data_out = 8'hBE;
                    16'hE225: data_out = 8'hBD;
                    16'hE226: data_out = 8'hBC;
                    16'hE227: data_out = 8'hBB;
                    16'hE228: data_out = 8'hBA;
                    16'hE229: data_out = 8'hB9;
                    16'hE22A: data_out = 8'hB8;
                    16'hE22B: data_out = 8'hB7;
                    16'hE22C: data_out = 8'hB6;
                    16'hE22D: data_out = 8'hB5;
                    16'hE22E: data_out = 8'hB4;
                    16'hE22F: data_out = 8'hB3;
                    16'hE230: data_out = 8'hB2;
                    16'hE231: data_out = 8'hB1;
                    16'hE232: data_out = 8'hB0;
                    16'hE233: data_out = 8'hAF;
                    16'hE234: data_out = 8'hAE;
                    16'hE235: data_out = 8'hAD;
                    16'hE236: data_out = 8'hAC;
                    16'hE237: data_out = 8'hAB;
                    16'hE238: data_out = 8'hAA;
                    16'hE239: data_out = 8'hA9;
                    16'hE23A: data_out = 8'hA8;
                    16'hE23B: data_out = 8'hA7;
                    16'hE23C: data_out = 8'hA6;
                    16'hE23D: data_out = 8'hA5;
                    16'hE23E: data_out = 8'hA4;
                    16'hE23F: data_out = 8'hA3;
                    16'hE240: data_out = 8'hA2;
                    16'hE241: data_out = 8'hA1;
                    16'hE242: data_out = 8'hA0;
                    16'hE243: data_out = 8'h9F;
                    16'hE244: data_out = 8'h9E;
                    16'hE245: data_out = 8'h9D;
                    16'hE246: data_out = 8'h9C;
                    16'hE247: data_out = 8'h9B;
                    16'hE248: data_out = 8'h9A;
                    16'hE249: data_out = 8'h99;
                    16'hE24A: data_out = 8'h98;
                    16'hE24B: data_out = 8'h97;
                    16'hE24C: data_out = 8'h96;
                    16'hE24D: data_out = 8'h95;
                    16'hE24E: data_out = 8'h94;
                    16'hE24F: data_out = 8'h93;
                    16'hE250: data_out = 8'h92;
                    16'hE251: data_out = 8'h91;
                    16'hE252: data_out = 8'h90;
                    16'hE253: data_out = 8'h8F;
                    16'hE254: data_out = 8'h8E;
                    16'hE255: data_out = 8'h8D;
                    16'hE256: data_out = 8'h8C;
                    16'hE257: data_out = 8'h8B;
                    16'hE258: data_out = 8'h8A;
                    16'hE259: data_out = 8'h89;
                    16'hE25A: data_out = 8'h88;
                    16'hE25B: data_out = 8'h87;
                    16'hE25C: data_out = 8'h86;
                    16'hE25D: data_out = 8'h85;
                    16'hE25E: data_out = 8'h84;
                    16'hE25F: data_out = 8'h83;
                    16'hE260: data_out = 8'h82;
                    16'hE261: data_out = 8'h81;
                    16'hE262: data_out = 8'h0;
                    16'hE263: data_out = 8'h1;
                    16'hE264: data_out = 8'h2;
                    16'hE265: data_out = 8'h3;
                    16'hE266: data_out = 8'h4;
                    16'hE267: data_out = 8'h5;
                    16'hE268: data_out = 8'h6;
                    16'hE269: data_out = 8'h7;
                    16'hE26A: data_out = 8'h8;
                    16'hE26B: data_out = 8'h9;
                    16'hE26C: data_out = 8'hA;
                    16'hE26D: data_out = 8'hB;
                    16'hE26E: data_out = 8'hC;
                    16'hE26F: data_out = 8'hD;
                    16'hE270: data_out = 8'hE;
                    16'hE271: data_out = 8'hF;
                    16'hE272: data_out = 8'h10;
                    16'hE273: data_out = 8'h11;
                    16'hE274: data_out = 8'h12;
                    16'hE275: data_out = 8'h13;
                    16'hE276: data_out = 8'h14;
                    16'hE277: data_out = 8'h15;
                    16'hE278: data_out = 8'h16;
                    16'hE279: data_out = 8'h17;
                    16'hE27A: data_out = 8'h18;
                    16'hE27B: data_out = 8'h19;
                    16'hE27C: data_out = 8'h1A;
                    16'hE27D: data_out = 8'h1B;
                    16'hE27E: data_out = 8'h1C;
                    16'hE27F: data_out = 8'h1D;
                    16'hE280: data_out = 8'hE2;
                    16'hE281: data_out = 8'hE3;
                    16'hE282: data_out = 8'hE4;
                    16'hE283: data_out = 8'hE5;
                    16'hE284: data_out = 8'hE6;
                    16'hE285: data_out = 8'hE7;
                    16'hE286: data_out = 8'hE8;
                    16'hE287: data_out = 8'hE9;
                    16'hE288: data_out = 8'hEA;
                    16'hE289: data_out = 8'hEB;
                    16'hE28A: data_out = 8'hEC;
                    16'hE28B: data_out = 8'hED;
                    16'hE28C: data_out = 8'hEE;
                    16'hE28D: data_out = 8'hEF;
                    16'hE28E: data_out = 8'hF0;
                    16'hE28F: data_out = 8'hF1;
                    16'hE290: data_out = 8'hF2;
                    16'hE291: data_out = 8'hF3;
                    16'hE292: data_out = 8'hF4;
                    16'hE293: data_out = 8'hF5;
                    16'hE294: data_out = 8'hF6;
                    16'hE295: data_out = 8'hF7;
                    16'hE296: data_out = 8'hF8;
                    16'hE297: data_out = 8'hF9;
                    16'hE298: data_out = 8'hFA;
                    16'hE299: data_out = 8'hFB;
                    16'hE29A: data_out = 8'hFC;
                    16'hE29B: data_out = 8'hFD;
                    16'hE29C: data_out = 8'hFE;
                    16'hE29D: data_out = 8'hFF;
                    16'hE29E: data_out = 8'h80;
                    16'hE29F: data_out = 8'h81;
                    16'hE2A0: data_out = 8'h82;
                    16'hE2A1: data_out = 8'h83;
                    16'hE2A2: data_out = 8'h84;
                    16'hE2A3: data_out = 8'h85;
                    16'hE2A4: data_out = 8'h86;
                    16'hE2A5: data_out = 8'h87;
                    16'hE2A6: data_out = 8'h88;
                    16'hE2A7: data_out = 8'h89;
                    16'hE2A8: data_out = 8'h8A;
                    16'hE2A9: data_out = 8'h8B;
                    16'hE2AA: data_out = 8'h8C;
                    16'hE2AB: data_out = 8'h8D;
                    16'hE2AC: data_out = 8'h8E;
                    16'hE2AD: data_out = 8'h8F;
                    16'hE2AE: data_out = 8'h90;
                    16'hE2AF: data_out = 8'h91;
                    16'hE2B0: data_out = 8'h92;
                    16'hE2B1: data_out = 8'h93;
                    16'hE2B2: data_out = 8'h94;
                    16'hE2B3: data_out = 8'h95;
                    16'hE2B4: data_out = 8'h96;
                    16'hE2B5: data_out = 8'h97;
                    16'hE2B6: data_out = 8'h98;
                    16'hE2B7: data_out = 8'h99;
                    16'hE2B8: data_out = 8'h9A;
                    16'hE2B9: data_out = 8'h9B;
                    16'hE2BA: data_out = 8'h9C;
                    16'hE2BB: data_out = 8'h9D;
                    16'hE2BC: data_out = 8'h9E;
                    16'hE2BD: data_out = 8'h9F;
                    16'hE2BE: data_out = 8'hA0;
                    16'hE2BF: data_out = 8'hA1;
                    16'hE2C0: data_out = 8'hA2;
                    16'hE2C1: data_out = 8'hA3;
                    16'hE2C2: data_out = 8'hA4;
                    16'hE2C3: data_out = 8'hA5;
                    16'hE2C4: data_out = 8'hA6;
                    16'hE2C5: data_out = 8'hA7;
                    16'hE2C6: data_out = 8'hA8;
                    16'hE2C7: data_out = 8'hA9;
                    16'hE2C8: data_out = 8'hAA;
                    16'hE2C9: data_out = 8'hAB;
                    16'hE2CA: data_out = 8'hAC;
                    16'hE2CB: data_out = 8'hAD;
                    16'hE2CC: data_out = 8'hAE;
                    16'hE2CD: data_out = 8'hAF;
                    16'hE2CE: data_out = 8'hB0;
                    16'hE2CF: data_out = 8'hB1;
                    16'hE2D0: data_out = 8'hB2;
                    16'hE2D1: data_out = 8'hB3;
                    16'hE2D2: data_out = 8'hB4;
                    16'hE2D3: data_out = 8'hB5;
                    16'hE2D4: data_out = 8'hB6;
                    16'hE2D5: data_out = 8'hB7;
                    16'hE2D6: data_out = 8'hB8;
                    16'hE2D7: data_out = 8'hB9;
                    16'hE2D8: data_out = 8'hBA;
                    16'hE2D9: data_out = 8'hBB;
                    16'hE2DA: data_out = 8'hBC;
                    16'hE2DB: data_out = 8'hBD;
                    16'hE2DC: data_out = 8'hBE;
                    16'hE2DD: data_out = 8'hBF;
                    16'hE2DE: data_out = 8'hC0;
                    16'hE2DF: data_out = 8'hC1;
                    16'hE2E0: data_out = 8'hC2;
                    16'hE2E1: data_out = 8'hC3;
                    16'hE2E2: data_out = 8'hC4;
                    16'hE2E3: data_out = 8'hC5;
                    16'hE2E4: data_out = 8'hC6;
                    16'hE2E5: data_out = 8'hC7;
                    16'hE2E6: data_out = 8'hC8;
                    16'hE2E7: data_out = 8'hC9;
                    16'hE2E8: data_out = 8'hCA;
                    16'hE2E9: data_out = 8'hCB;
                    16'hE2EA: data_out = 8'hCC;
                    16'hE2EB: data_out = 8'hCD;
                    16'hE2EC: data_out = 8'hCE;
                    16'hE2ED: data_out = 8'hCF;
                    16'hE2EE: data_out = 8'hD0;
                    16'hE2EF: data_out = 8'hD1;
                    16'hE2F0: data_out = 8'hD2;
                    16'hE2F1: data_out = 8'hD3;
                    16'hE2F2: data_out = 8'hD4;
                    16'hE2F3: data_out = 8'hD5;
                    16'hE2F4: data_out = 8'hD6;
                    16'hE2F5: data_out = 8'hD7;
                    16'hE2F6: data_out = 8'hD8;
                    16'hE2F7: data_out = 8'hD9;
                    16'hE2F8: data_out = 8'hDA;
                    16'hE2F9: data_out = 8'hDB;
                    16'hE2FA: data_out = 8'hDC;
                    16'hE2FB: data_out = 8'hDD;
                    16'hE2FC: data_out = 8'hDE;
                    16'hE2FD: data_out = 8'hDF;
                    16'hE2FE: data_out = 8'hE0;
                    16'hE2FF: data_out = 8'hE1;
                    16'hE300: data_out = 8'hE3;
                    16'hE301: data_out = 8'hE2;
                    16'hE302: data_out = 8'hE1;
                    16'hE303: data_out = 8'hE0;
                    16'hE304: data_out = 8'hDF;
                    16'hE305: data_out = 8'hDE;
                    16'hE306: data_out = 8'hDD;
                    16'hE307: data_out = 8'hDC;
                    16'hE308: data_out = 8'hDB;
                    16'hE309: data_out = 8'hDA;
                    16'hE30A: data_out = 8'hD9;
                    16'hE30B: data_out = 8'hD8;
                    16'hE30C: data_out = 8'hD7;
                    16'hE30D: data_out = 8'hD6;
                    16'hE30E: data_out = 8'hD5;
                    16'hE30F: data_out = 8'hD4;
                    16'hE310: data_out = 8'hD3;
                    16'hE311: data_out = 8'hD2;
                    16'hE312: data_out = 8'hD1;
                    16'hE313: data_out = 8'hD0;
                    16'hE314: data_out = 8'hCF;
                    16'hE315: data_out = 8'hCE;
                    16'hE316: data_out = 8'hCD;
                    16'hE317: data_out = 8'hCC;
                    16'hE318: data_out = 8'hCB;
                    16'hE319: data_out = 8'hCA;
                    16'hE31A: data_out = 8'hC9;
                    16'hE31B: data_out = 8'hC8;
                    16'hE31C: data_out = 8'hC7;
                    16'hE31D: data_out = 8'hC6;
                    16'hE31E: data_out = 8'hC5;
                    16'hE31F: data_out = 8'hC4;
                    16'hE320: data_out = 8'hC3;
                    16'hE321: data_out = 8'hC2;
                    16'hE322: data_out = 8'hC1;
                    16'hE323: data_out = 8'hC0;
                    16'hE324: data_out = 8'hBF;
                    16'hE325: data_out = 8'hBE;
                    16'hE326: data_out = 8'hBD;
                    16'hE327: data_out = 8'hBC;
                    16'hE328: data_out = 8'hBB;
                    16'hE329: data_out = 8'hBA;
                    16'hE32A: data_out = 8'hB9;
                    16'hE32B: data_out = 8'hB8;
                    16'hE32C: data_out = 8'hB7;
                    16'hE32D: data_out = 8'hB6;
                    16'hE32E: data_out = 8'hB5;
                    16'hE32F: data_out = 8'hB4;
                    16'hE330: data_out = 8'hB3;
                    16'hE331: data_out = 8'hB2;
                    16'hE332: data_out = 8'hB1;
                    16'hE333: data_out = 8'hB0;
                    16'hE334: data_out = 8'hAF;
                    16'hE335: data_out = 8'hAE;
                    16'hE336: data_out = 8'hAD;
                    16'hE337: data_out = 8'hAC;
                    16'hE338: data_out = 8'hAB;
                    16'hE339: data_out = 8'hAA;
                    16'hE33A: data_out = 8'hA9;
                    16'hE33B: data_out = 8'hA8;
                    16'hE33C: data_out = 8'hA7;
                    16'hE33D: data_out = 8'hA6;
                    16'hE33E: data_out = 8'hA5;
                    16'hE33F: data_out = 8'hA4;
                    16'hE340: data_out = 8'hA3;
                    16'hE341: data_out = 8'hA2;
                    16'hE342: data_out = 8'hA1;
                    16'hE343: data_out = 8'hA0;
                    16'hE344: data_out = 8'h9F;
                    16'hE345: data_out = 8'h9E;
                    16'hE346: data_out = 8'h9D;
                    16'hE347: data_out = 8'h9C;
                    16'hE348: data_out = 8'h9B;
                    16'hE349: data_out = 8'h9A;
                    16'hE34A: data_out = 8'h99;
                    16'hE34B: data_out = 8'h98;
                    16'hE34C: data_out = 8'h97;
                    16'hE34D: data_out = 8'h96;
                    16'hE34E: data_out = 8'h95;
                    16'hE34F: data_out = 8'h94;
                    16'hE350: data_out = 8'h93;
                    16'hE351: data_out = 8'h92;
                    16'hE352: data_out = 8'h91;
                    16'hE353: data_out = 8'h90;
                    16'hE354: data_out = 8'h8F;
                    16'hE355: data_out = 8'h8E;
                    16'hE356: data_out = 8'h8D;
                    16'hE357: data_out = 8'h8C;
                    16'hE358: data_out = 8'h8B;
                    16'hE359: data_out = 8'h8A;
                    16'hE35A: data_out = 8'h89;
                    16'hE35B: data_out = 8'h88;
                    16'hE35C: data_out = 8'h87;
                    16'hE35D: data_out = 8'h86;
                    16'hE35E: data_out = 8'h85;
                    16'hE35F: data_out = 8'h84;
                    16'hE360: data_out = 8'h83;
                    16'hE361: data_out = 8'h82;
                    16'hE362: data_out = 8'h81;
                    16'hE363: data_out = 8'h0;
                    16'hE364: data_out = 8'h1;
                    16'hE365: data_out = 8'h2;
                    16'hE366: data_out = 8'h3;
                    16'hE367: data_out = 8'h4;
                    16'hE368: data_out = 8'h5;
                    16'hE369: data_out = 8'h6;
                    16'hE36A: data_out = 8'h7;
                    16'hE36B: data_out = 8'h8;
                    16'hE36C: data_out = 8'h9;
                    16'hE36D: data_out = 8'hA;
                    16'hE36E: data_out = 8'hB;
                    16'hE36F: data_out = 8'hC;
                    16'hE370: data_out = 8'hD;
                    16'hE371: data_out = 8'hE;
                    16'hE372: data_out = 8'hF;
                    16'hE373: data_out = 8'h10;
                    16'hE374: data_out = 8'h11;
                    16'hE375: data_out = 8'h12;
                    16'hE376: data_out = 8'h13;
                    16'hE377: data_out = 8'h14;
                    16'hE378: data_out = 8'h15;
                    16'hE379: data_out = 8'h16;
                    16'hE37A: data_out = 8'h17;
                    16'hE37B: data_out = 8'h18;
                    16'hE37C: data_out = 8'h19;
                    16'hE37D: data_out = 8'h1A;
                    16'hE37E: data_out = 8'h1B;
                    16'hE37F: data_out = 8'h1C;
                    16'hE380: data_out = 8'hE3;
                    16'hE381: data_out = 8'hE4;
                    16'hE382: data_out = 8'hE5;
                    16'hE383: data_out = 8'hE6;
                    16'hE384: data_out = 8'hE7;
                    16'hE385: data_out = 8'hE8;
                    16'hE386: data_out = 8'hE9;
                    16'hE387: data_out = 8'hEA;
                    16'hE388: data_out = 8'hEB;
                    16'hE389: data_out = 8'hEC;
                    16'hE38A: data_out = 8'hED;
                    16'hE38B: data_out = 8'hEE;
                    16'hE38C: data_out = 8'hEF;
                    16'hE38D: data_out = 8'hF0;
                    16'hE38E: data_out = 8'hF1;
                    16'hE38F: data_out = 8'hF2;
                    16'hE390: data_out = 8'hF3;
                    16'hE391: data_out = 8'hF4;
                    16'hE392: data_out = 8'hF5;
                    16'hE393: data_out = 8'hF6;
                    16'hE394: data_out = 8'hF7;
                    16'hE395: data_out = 8'hF8;
                    16'hE396: data_out = 8'hF9;
                    16'hE397: data_out = 8'hFA;
                    16'hE398: data_out = 8'hFB;
                    16'hE399: data_out = 8'hFC;
                    16'hE39A: data_out = 8'hFD;
                    16'hE39B: data_out = 8'hFE;
                    16'hE39C: data_out = 8'hFF;
                    16'hE39D: data_out = 8'h80;
                    16'hE39E: data_out = 8'h81;
                    16'hE39F: data_out = 8'h82;
                    16'hE3A0: data_out = 8'h83;
                    16'hE3A1: data_out = 8'h84;
                    16'hE3A2: data_out = 8'h85;
                    16'hE3A3: data_out = 8'h86;
                    16'hE3A4: data_out = 8'h87;
                    16'hE3A5: data_out = 8'h88;
                    16'hE3A6: data_out = 8'h89;
                    16'hE3A7: data_out = 8'h8A;
                    16'hE3A8: data_out = 8'h8B;
                    16'hE3A9: data_out = 8'h8C;
                    16'hE3AA: data_out = 8'h8D;
                    16'hE3AB: data_out = 8'h8E;
                    16'hE3AC: data_out = 8'h8F;
                    16'hE3AD: data_out = 8'h90;
                    16'hE3AE: data_out = 8'h91;
                    16'hE3AF: data_out = 8'h92;
                    16'hE3B0: data_out = 8'h93;
                    16'hE3B1: data_out = 8'h94;
                    16'hE3B2: data_out = 8'h95;
                    16'hE3B3: data_out = 8'h96;
                    16'hE3B4: data_out = 8'h97;
                    16'hE3B5: data_out = 8'h98;
                    16'hE3B6: data_out = 8'h99;
                    16'hE3B7: data_out = 8'h9A;
                    16'hE3B8: data_out = 8'h9B;
                    16'hE3B9: data_out = 8'h9C;
                    16'hE3BA: data_out = 8'h9D;
                    16'hE3BB: data_out = 8'h9E;
                    16'hE3BC: data_out = 8'h9F;
                    16'hE3BD: data_out = 8'hA0;
                    16'hE3BE: data_out = 8'hA1;
                    16'hE3BF: data_out = 8'hA2;
                    16'hE3C0: data_out = 8'hA3;
                    16'hE3C1: data_out = 8'hA4;
                    16'hE3C2: data_out = 8'hA5;
                    16'hE3C3: data_out = 8'hA6;
                    16'hE3C4: data_out = 8'hA7;
                    16'hE3C5: data_out = 8'hA8;
                    16'hE3C6: data_out = 8'hA9;
                    16'hE3C7: data_out = 8'hAA;
                    16'hE3C8: data_out = 8'hAB;
                    16'hE3C9: data_out = 8'hAC;
                    16'hE3CA: data_out = 8'hAD;
                    16'hE3CB: data_out = 8'hAE;
                    16'hE3CC: data_out = 8'hAF;
                    16'hE3CD: data_out = 8'hB0;
                    16'hE3CE: data_out = 8'hB1;
                    16'hE3CF: data_out = 8'hB2;
                    16'hE3D0: data_out = 8'hB3;
                    16'hE3D1: data_out = 8'hB4;
                    16'hE3D2: data_out = 8'hB5;
                    16'hE3D3: data_out = 8'hB6;
                    16'hE3D4: data_out = 8'hB7;
                    16'hE3D5: data_out = 8'hB8;
                    16'hE3D6: data_out = 8'hB9;
                    16'hE3D7: data_out = 8'hBA;
                    16'hE3D8: data_out = 8'hBB;
                    16'hE3D9: data_out = 8'hBC;
                    16'hE3DA: data_out = 8'hBD;
                    16'hE3DB: data_out = 8'hBE;
                    16'hE3DC: data_out = 8'hBF;
                    16'hE3DD: data_out = 8'hC0;
                    16'hE3DE: data_out = 8'hC1;
                    16'hE3DF: data_out = 8'hC2;
                    16'hE3E0: data_out = 8'hC3;
                    16'hE3E1: data_out = 8'hC4;
                    16'hE3E2: data_out = 8'hC5;
                    16'hE3E3: data_out = 8'hC6;
                    16'hE3E4: data_out = 8'hC7;
                    16'hE3E5: data_out = 8'hC8;
                    16'hE3E6: data_out = 8'hC9;
                    16'hE3E7: data_out = 8'hCA;
                    16'hE3E8: data_out = 8'hCB;
                    16'hE3E9: data_out = 8'hCC;
                    16'hE3EA: data_out = 8'hCD;
                    16'hE3EB: data_out = 8'hCE;
                    16'hE3EC: data_out = 8'hCF;
                    16'hE3ED: data_out = 8'hD0;
                    16'hE3EE: data_out = 8'hD1;
                    16'hE3EF: data_out = 8'hD2;
                    16'hE3F0: data_out = 8'hD3;
                    16'hE3F1: data_out = 8'hD4;
                    16'hE3F2: data_out = 8'hD5;
                    16'hE3F3: data_out = 8'hD6;
                    16'hE3F4: data_out = 8'hD7;
                    16'hE3F5: data_out = 8'hD8;
                    16'hE3F6: data_out = 8'hD9;
                    16'hE3F7: data_out = 8'hDA;
                    16'hE3F8: data_out = 8'hDB;
                    16'hE3F9: data_out = 8'hDC;
                    16'hE3FA: data_out = 8'hDD;
                    16'hE3FB: data_out = 8'hDE;
                    16'hE3FC: data_out = 8'hDF;
                    16'hE3FD: data_out = 8'hE0;
                    16'hE3FE: data_out = 8'hE1;
                    16'hE3FF: data_out = 8'hE2;
                    16'hE400: data_out = 8'hE4;
                    16'hE401: data_out = 8'hE3;
                    16'hE402: data_out = 8'hE2;
                    16'hE403: data_out = 8'hE1;
                    16'hE404: data_out = 8'hE0;
                    16'hE405: data_out = 8'hDF;
                    16'hE406: data_out = 8'hDE;
                    16'hE407: data_out = 8'hDD;
                    16'hE408: data_out = 8'hDC;
                    16'hE409: data_out = 8'hDB;
                    16'hE40A: data_out = 8'hDA;
                    16'hE40B: data_out = 8'hD9;
                    16'hE40C: data_out = 8'hD8;
                    16'hE40D: data_out = 8'hD7;
                    16'hE40E: data_out = 8'hD6;
                    16'hE40F: data_out = 8'hD5;
                    16'hE410: data_out = 8'hD4;
                    16'hE411: data_out = 8'hD3;
                    16'hE412: data_out = 8'hD2;
                    16'hE413: data_out = 8'hD1;
                    16'hE414: data_out = 8'hD0;
                    16'hE415: data_out = 8'hCF;
                    16'hE416: data_out = 8'hCE;
                    16'hE417: data_out = 8'hCD;
                    16'hE418: data_out = 8'hCC;
                    16'hE419: data_out = 8'hCB;
                    16'hE41A: data_out = 8'hCA;
                    16'hE41B: data_out = 8'hC9;
                    16'hE41C: data_out = 8'hC8;
                    16'hE41D: data_out = 8'hC7;
                    16'hE41E: data_out = 8'hC6;
                    16'hE41F: data_out = 8'hC5;
                    16'hE420: data_out = 8'hC4;
                    16'hE421: data_out = 8'hC3;
                    16'hE422: data_out = 8'hC2;
                    16'hE423: data_out = 8'hC1;
                    16'hE424: data_out = 8'hC0;
                    16'hE425: data_out = 8'hBF;
                    16'hE426: data_out = 8'hBE;
                    16'hE427: data_out = 8'hBD;
                    16'hE428: data_out = 8'hBC;
                    16'hE429: data_out = 8'hBB;
                    16'hE42A: data_out = 8'hBA;
                    16'hE42B: data_out = 8'hB9;
                    16'hE42C: data_out = 8'hB8;
                    16'hE42D: data_out = 8'hB7;
                    16'hE42E: data_out = 8'hB6;
                    16'hE42F: data_out = 8'hB5;
                    16'hE430: data_out = 8'hB4;
                    16'hE431: data_out = 8'hB3;
                    16'hE432: data_out = 8'hB2;
                    16'hE433: data_out = 8'hB1;
                    16'hE434: data_out = 8'hB0;
                    16'hE435: data_out = 8'hAF;
                    16'hE436: data_out = 8'hAE;
                    16'hE437: data_out = 8'hAD;
                    16'hE438: data_out = 8'hAC;
                    16'hE439: data_out = 8'hAB;
                    16'hE43A: data_out = 8'hAA;
                    16'hE43B: data_out = 8'hA9;
                    16'hE43C: data_out = 8'hA8;
                    16'hE43D: data_out = 8'hA7;
                    16'hE43E: data_out = 8'hA6;
                    16'hE43F: data_out = 8'hA5;
                    16'hE440: data_out = 8'hA4;
                    16'hE441: data_out = 8'hA3;
                    16'hE442: data_out = 8'hA2;
                    16'hE443: data_out = 8'hA1;
                    16'hE444: data_out = 8'hA0;
                    16'hE445: data_out = 8'h9F;
                    16'hE446: data_out = 8'h9E;
                    16'hE447: data_out = 8'h9D;
                    16'hE448: data_out = 8'h9C;
                    16'hE449: data_out = 8'h9B;
                    16'hE44A: data_out = 8'h9A;
                    16'hE44B: data_out = 8'h99;
                    16'hE44C: data_out = 8'h98;
                    16'hE44D: data_out = 8'h97;
                    16'hE44E: data_out = 8'h96;
                    16'hE44F: data_out = 8'h95;
                    16'hE450: data_out = 8'h94;
                    16'hE451: data_out = 8'h93;
                    16'hE452: data_out = 8'h92;
                    16'hE453: data_out = 8'h91;
                    16'hE454: data_out = 8'h90;
                    16'hE455: data_out = 8'h8F;
                    16'hE456: data_out = 8'h8E;
                    16'hE457: data_out = 8'h8D;
                    16'hE458: data_out = 8'h8C;
                    16'hE459: data_out = 8'h8B;
                    16'hE45A: data_out = 8'h8A;
                    16'hE45B: data_out = 8'h89;
                    16'hE45C: data_out = 8'h88;
                    16'hE45D: data_out = 8'h87;
                    16'hE45E: data_out = 8'h86;
                    16'hE45F: data_out = 8'h85;
                    16'hE460: data_out = 8'h84;
                    16'hE461: data_out = 8'h83;
                    16'hE462: data_out = 8'h82;
                    16'hE463: data_out = 8'h81;
                    16'hE464: data_out = 8'h0;
                    16'hE465: data_out = 8'h1;
                    16'hE466: data_out = 8'h2;
                    16'hE467: data_out = 8'h3;
                    16'hE468: data_out = 8'h4;
                    16'hE469: data_out = 8'h5;
                    16'hE46A: data_out = 8'h6;
                    16'hE46B: data_out = 8'h7;
                    16'hE46C: data_out = 8'h8;
                    16'hE46D: data_out = 8'h9;
                    16'hE46E: data_out = 8'hA;
                    16'hE46F: data_out = 8'hB;
                    16'hE470: data_out = 8'hC;
                    16'hE471: data_out = 8'hD;
                    16'hE472: data_out = 8'hE;
                    16'hE473: data_out = 8'hF;
                    16'hE474: data_out = 8'h10;
                    16'hE475: data_out = 8'h11;
                    16'hE476: data_out = 8'h12;
                    16'hE477: data_out = 8'h13;
                    16'hE478: data_out = 8'h14;
                    16'hE479: data_out = 8'h15;
                    16'hE47A: data_out = 8'h16;
                    16'hE47B: data_out = 8'h17;
                    16'hE47C: data_out = 8'h18;
                    16'hE47D: data_out = 8'h19;
                    16'hE47E: data_out = 8'h1A;
                    16'hE47F: data_out = 8'h1B;
                    16'hE480: data_out = 8'hE4;
                    16'hE481: data_out = 8'hE5;
                    16'hE482: data_out = 8'hE6;
                    16'hE483: data_out = 8'hE7;
                    16'hE484: data_out = 8'hE8;
                    16'hE485: data_out = 8'hE9;
                    16'hE486: data_out = 8'hEA;
                    16'hE487: data_out = 8'hEB;
                    16'hE488: data_out = 8'hEC;
                    16'hE489: data_out = 8'hED;
                    16'hE48A: data_out = 8'hEE;
                    16'hE48B: data_out = 8'hEF;
                    16'hE48C: data_out = 8'hF0;
                    16'hE48D: data_out = 8'hF1;
                    16'hE48E: data_out = 8'hF2;
                    16'hE48F: data_out = 8'hF3;
                    16'hE490: data_out = 8'hF4;
                    16'hE491: data_out = 8'hF5;
                    16'hE492: data_out = 8'hF6;
                    16'hE493: data_out = 8'hF7;
                    16'hE494: data_out = 8'hF8;
                    16'hE495: data_out = 8'hF9;
                    16'hE496: data_out = 8'hFA;
                    16'hE497: data_out = 8'hFB;
                    16'hE498: data_out = 8'hFC;
                    16'hE499: data_out = 8'hFD;
                    16'hE49A: data_out = 8'hFE;
                    16'hE49B: data_out = 8'hFF;
                    16'hE49C: data_out = 8'h80;
                    16'hE49D: data_out = 8'h81;
                    16'hE49E: data_out = 8'h82;
                    16'hE49F: data_out = 8'h83;
                    16'hE4A0: data_out = 8'h84;
                    16'hE4A1: data_out = 8'h85;
                    16'hE4A2: data_out = 8'h86;
                    16'hE4A3: data_out = 8'h87;
                    16'hE4A4: data_out = 8'h88;
                    16'hE4A5: data_out = 8'h89;
                    16'hE4A6: data_out = 8'h8A;
                    16'hE4A7: data_out = 8'h8B;
                    16'hE4A8: data_out = 8'h8C;
                    16'hE4A9: data_out = 8'h8D;
                    16'hE4AA: data_out = 8'h8E;
                    16'hE4AB: data_out = 8'h8F;
                    16'hE4AC: data_out = 8'h90;
                    16'hE4AD: data_out = 8'h91;
                    16'hE4AE: data_out = 8'h92;
                    16'hE4AF: data_out = 8'h93;
                    16'hE4B0: data_out = 8'h94;
                    16'hE4B1: data_out = 8'h95;
                    16'hE4B2: data_out = 8'h96;
                    16'hE4B3: data_out = 8'h97;
                    16'hE4B4: data_out = 8'h98;
                    16'hE4B5: data_out = 8'h99;
                    16'hE4B6: data_out = 8'h9A;
                    16'hE4B7: data_out = 8'h9B;
                    16'hE4B8: data_out = 8'h9C;
                    16'hE4B9: data_out = 8'h9D;
                    16'hE4BA: data_out = 8'h9E;
                    16'hE4BB: data_out = 8'h9F;
                    16'hE4BC: data_out = 8'hA0;
                    16'hE4BD: data_out = 8'hA1;
                    16'hE4BE: data_out = 8'hA2;
                    16'hE4BF: data_out = 8'hA3;
                    16'hE4C0: data_out = 8'hA4;
                    16'hE4C1: data_out = 8'hA5;
                    16'hE4C2: data_out = 8'hA6;
                    16'hE4C3: data_out = 8'hA7;
                    16'hE4C4: data_out = 8'hA8;
                    16'hE4C5: data_out = 8'hA9;
                    16'hE4C6: data_out = 8'hAA;
                    16'hE4C7: data_out = 8'hAB;
                    16'hE4C8: data_out = 8'hAC;
                    16'hE4C9: data_out = 8'hAD;
                    16'hE4CA: data_out = 8'hAE;
                    16'hE4CB: data_out = 8'hAF;
                    16'hE4CC: data_out = 8'hB0;
                    16'hE4CD: data_out = 8'hB1;
                    16'hE4CE: data_out = 8'hB2;
                    16'hE4CF: data_out = 8'hB3;
                    16'hE4D0: data_out = 8'hB4;
                    16'hE4D1: data_out = 8'hB5;
                    16'hE4D2: data_out = 8'hB6;
                    16'hE4D3: data_out = 8'hB7;
                    16'hE4D4: data_out = 8'hB8;
                    16'hE4D5: data_out = 8'hB9;
                    16'hE4D6: data_out = 8'hBA;
                    16'hE4D7: data_out = 8'hBB;
                    16'hE4D8: data_out = 8'hBC;
                    16'hE4D9: data_out = 8'hBD;
                    16'hE4DA: data_out = 8'hBE;
                    16'hE4DB: data_out = 8'hBF;
                    16'hE4DC: data_out = 8'hC0;
                    16'hE4DD: data_out = 8'hC1;
                    16'hE4DE: data_out = 8'hC2;
                    16'hE4DF: data_out = 8'hC3;
                    16'hE4E0: data_out = 8'hC4;
                    16'hE4E1: data_out = 8'hC5;
                    16'hE4E2: data_out = 8'hC6;
                    16'hE4E3: data_out = 8'hC7;
                    16'hE4E4: data_out = 8'hC8;
                    16'hE4E5: data_out = 8'hC9;
                    16'hE4E6: data_out = 8'hCA;
                    16'hE4E7: data_out = 8'hCB;
                    16'hE4E8: data_out = 8'hCC;
                    16'hE4E9: data_out = 8'hCD;
                    16'hE4EA: data_out = 8'hCE;
                    16'hE4EB: data_out = 8'hCF;
                    16'hE4EC: data_out = 8'hD0;
                    16'hE4ED: data_out = 8'hD1;
                    16'hE4EE: data_out = 8'hD2;
                    16'hE4EF: data_out = 8'hD3;
                    16'hE4F0: data_out = 8'hD4;
                    16'hE4F1: data_out = 8'hD5;
                    16'hE4F2: data_out = 8'hD6;
                    16'hE4F3: data_out = 8'hD7;
                    16'hE4F4: data_out = 8'hD8;
                    16'hE4F5: data_out = 8'hD9;
                    16'hE4F6: data_out = 8'hDA;
                    16'hE4F7: data_out = 8'hDB;
                    16'hE4F8: data_out = 8'hDC;
                    16'hE4F9: data_out = 8'hDD;
                    16'hE4FA: data_out = 8'hDE;
                    16'hE4FB: data_out = 8'hDF;
                    16'hE4FC: data_out = 8'hE0;
                    16'hE4FD: data_out = 8'hE1;
                    16'hE4FE: data_out = 8'hE2;
                    16'hE4FF: data_out = 8'hE3;
                    16'hE500: data_out = 8'hE5;
                    16'hE501: data_out = 8'hE4;
                    16'hE502: data_out = 8'hE3;
                    16'hE503: data_out = 8'hE2;
                    16'hE504: data_out = 8'hE1;
                    16'hE505: data_out = 8'hE0;
                    16'hE506: data_out = 8'hDF;
                    16'hE507: data_out = 8'hDE;
                    16'hE508: data_out = 8'hDD;
                    16'hE509: data_out = 8'hDC;
                    16'hE50A: data_out = 8'hDB;
                    16'hE50B: data_out = 8'hDA;
                    16'hE50C: data_out = 8'hD9;
                    16'hE50D: data_out = 8'hD8;
                    16'hE50E: data_out = 8'hD7;
                    16'hE50F: data_out = 8'hD6;
                    16'hE510: data_out = 8'hD5;
                    16'hE511: data_out = 8'hD4;
                    16'hE512: data_out = 8'hD3;
                    16'hE513: data_out = 8'hD2;
                    16'hE514: data_out = 8'hD1;
                    16'hE515: data_out = 8'hD0;
                    16'hE516: data_out = 8'hCF;
                    16'hE517: data_out = 8'hCE;
                    16'hE518: data_out = 8'hCD;
                    16'hE519: data_out = 8'hCC;
                    16'hE51A: data_out = 8'hCB;
                    16'hE51B: data_out = 8'hCA;
                    16'hE51C: data_out = 8'hC9;
                    16'hE51D: data_out = 8'hC8;
                    16'hE51E: data_out = 8'hC7;
                    16'hE51F: data_out = 8'hC6;
                    16'hE520: data_out = 8'hC5;
                    16'hE521: data_out = 8'hC4;
                    16'hE522: data_out = 8'hC3;
                    16'hE523: data_out = 8'hC2;
                    16'hE524: data_out = 8'hC1;
                    16'hE525: data_out = 8'hC0;
                    16'hE526: data_out = 8'hBF;
                    16'hE527: data_out = 8'hBE;
                    16'hE528: data_out = 8'hBD;
                    16'hE529: data_out = 8'hBC;
                    16'hE52A: data_out = 8'hBB;
                    16'hE52B: data_out = 8'hBA;
                    16'hE52C: data_out = 8'hB9;
                    16'hE52D: data_out = 8'hB8;
                    16'hE52E: data_out = 8'hB7;
                    16'hE52F: data_out = 8'hB6;
                    16'hE530: data_out = 8'hB5;
                    16'hE531: data_out = 8'hB4;
                    16'hE532: data_out = 8'hB3;
                    16'hE533: data_out = 8'hB2;
                    16'hE534: data_out = 8'hB1;
                    16'hE535: data_out = 8'hB0;
                    16'hE536: data_out = 8'hAF;
                    16'hE537: data_out = 8'hAE;
                    16'hE538: data_out = 8'hAD;
                    16'hE539: data_out = 8'hAC;
                    16'hE53A: data_out = 8'hAB;
                    16'hE53B: data_out = 8'hAA;
                    16'hE53C: data_out = 8'hA9;
                    16'hE53D: data_out = 8'hA8;
                    16'hE53E: data_out = 8'hA7;
                    16'hE53F: data_out = 8'hA6;
                    16'hE540: data_out = 8'hA5;
                    16'hE541: data_out = 8'hA4;
                    16'hE542: data_out = 8'hA3;
                    16'hE543: data_out = 8'hA2;
                    16'hE544: data_out = 8'hA1;
                    16'hE545: data_out = 8'hA0;
                    16'hE546: data_out = 8'h9F;
                    16'hE547: data_out = 8'h9E;
                    16'hE548: data_out = 8'h9D;
                    16'hE549: data_out = 8'h9C;
                    16'hE54A: data_out = 8'h9B;
                    16'hE54B: data_out = 8'h9A;
                    16'hE54C: data_out = 8'h99;
                    16'hE54D: data_out = 8'h98;
                    16'hE54E: data_out = 8'h97;
                    16'hE54F: data_out = 8'h96;
                    16'hE550: data_out = 8'h95;
                    16'hE551: data_out = 8'h94;
                    16'hE552: data_out = 8'h93;
                    16'hE553: data_out = 8'h92;
                    16'hE554: data_out = 8'h91;
                    16'hE555: data_out = 8'h90;
                    16'hE556: data_out = 8'h8F;
                    16'hE557: data_out = 8'h8E;
                    16'hE558: data_out = 8'h8D;
                    16'hE559: data_out = 8'h8C;
                    16'hE55A: data_out = 8'h8B;
                    16'hE55B: data_out = 8'h8A;
                    16'hE55C: data_out = 8'h89;
                    16'hE55D: data_out = 8'h88;
                    16'hE55E: data_out = 8'h87;
                    16'hE55F: data_out = 8'h86;
                    16'hE560: data_out = 8'h85;
                    16'hE561: data_out = 8'h84;
                    16'hE562: data_out = 8'h83;
                    16'hE563: data_out = 8'h82;
                    16'hE564: data_out = 8'h81;
                    16'hE565: data_out = 8'h0;
                    16'hE566: data_out = 8'h1;
                    16'hE567: data_out = 8'h2;
                    16'hE568: data_out = 8'h3;
                    16'hE569: data_out = 8'h4;
                    16'hE56A: data_out = 8'h5;
                    16'hE56B: data_out = 8'h6;
                    16'hE56C: data_out = 8'h7;
                    16'hE56D: data_out = 8'h8;
                    16'hE56E: data_out = 8'h9;
                    16'hE56F: data_out = 8'hA;
                    16'hE570: data_out = 8'hB;
                    16'hE571: data_out = 8'hC;
                    16'hE572: data_out = 8'hD;
                    16'hE573: data_out = 8'hE;
                    16'hE574: data_out = 8'hF;
                    16'hE575: data_out = 8'h10;
                    16'hE576: data_out = 8'h11;
                    16'hE577: data_out = 8'h12;
                    16'hE578: data_out = 8'h13;
                    16'hE579: data_out = 8'h14;
                    16'hE57A: data_out = 8'h15;
                    16'hE57B: data_out = 8'h16;
                    16'hE57C: data_out = 8'h17;
                    16'hE57D: data_out = 8'h18;
                    16'hE57E: data_out = 8'h19;
                    16'hE57F: data_out = 8'h1A;
                    16'hE580: data_out = 8'hE5;
                    16'hE581: data_out = 8'hE6;
                    16'hE582: data_out = 8'hE7;
                    16'hE583: data_out = 8'hE8;
                    16'hE584: data_out = 8'hE9;
                    16'hE585: data_out = 8'hEA;
                    16'hE586: data_out = 8'hEB;
                    16'hE587: data_out = 8'hEC;
                    16'hE588: data_out = 8'hED;
                    16'hE589: data_out = 8'hEE;
                    16'hE58A: data_out = 8'hEF;
                    16'hE58B: data_out = 8'hF0;
                    16'hE58C: data_out = 8'hF1;
                    16'hE58D: data_out = 8'hF2;
                    16'hE58E: data_out = 8'hF3;
                    16'hE58F: data_out = 8'hF4;
                    16'hE590: data_out = 8'hF5;
                    16'hE591: data_out = 8'hF6;
                    16'hE592: data_out = 8'hF7;
                    16'hE593: data_out = 8'hF8;
                    16'hE594: data_out = 8'hF9;
                    16'hE595: data_out = 8'hFA;
                    16'hE596: data_out = 8'hFB;
                    16'hE597: data_out = 8'hFC;
                    16'hE598: data_out = 8'hFD;
                    16'hE599: data_out = 8'hFE;
                    16'hE59A: data_out = 8'hFF;
                    16'hE59B: data_out = 8'h80;
                    16'hE59C: data_out = 8'h81;
                    16'hE59D: data_out = 8'h82;
                    16'hE59E: data_out = 8'h83;
                    16'hE59F: data_out = 8'h84;
                    16'hE5A0: data_out = 8'h85;
                    16'hE5A1: data_out = 8'h86;
                    16'hE5A2: data_out = 8'h87;
                    16'hE5A3: data_out = 8'h88;
                    16'hE5A4: data_out = 8'h89;
                    16'hE5A5: data_out = 8'h8A;
                    16'hE5A6: data_out = 8'h8B;
                    16'hE5A7: data_out = 8'h8C;
                    16'hE5A8: data_out = 8'h8D;
                    16'hE5A9: data_out = 8'h8E;
                    16'hE5AA: data_out = 8'h8F;
                    16'hE5AB: data_out = 8'h90;
                    16'hE5AC: data_out = 8'h91;
                    16'hE5AD: data_out = 8'h92;
                    16'hE5AE: data_out = 8'h93;
                    16'hE5AF: data_out = 8'h94;
                    16'hE5B0: data_out = 8'h95;
                    16'hE5B1: data_out = 8'h96;
                    16'hE5B2: data_out = 8'h97;
                    16'hE5B3: data_out = 8'h98;
                    16'hE5B4: data_out = 8'h99;
                    16'hE5B5: data_out = 8'h9A;
                    16'hE5B6: data_out = 8'h9B;
                    16'hE5B7: data_out = 8'h9C;
                    16'hE5B8: data_out = 8'h9D;
                    16'hE5B9: data_out = 8'h9E;
                    16'hE5BA: data_out = 8'h9F;
                    16'hE5BB: data_out = 8'hA0;
                    16'hE5BC: data_out = 8'hA1;
                    16'hE5BD: data_out = 8'hA2;
                    16'hE5BE: data_out = 8'hA3;
                    16'hE5BF: data_out = 8'hA4;
                    16'hE5C0: data_out = 8'hA5;
                    16'hE5C1: data_out = 8'hA6;
                    16'hE5C2: data_out = 8'hA7;
                    16'hE5C3: data_out = 8'hA8;
                    16'hE5C4: data_out = 8'hA9;
                    16'hE5C5: data_out = 8'hAA;
                    16'hE5C6: data_out = 8'hAB;
                    16'hE5C7: data_out = 8'hAC;
                    16'hE5C8: data_out = 8'hAD;
                    16'hE5C9: data_out = 8'hAE;
                    16'hE5CA: data_out = 8'hAF;
                    16'hE5CB: data_out = 8'hB0;
                    16'hE5CC: data_out = 8'hB1;
                    16'hE5CD: data_out = 8'hB2;
                    16'hE5CE: data_out = 8'hB3;
                    16'hE5CF: data_out = 8'hB4;
                    16'hE5D0: data_out = 8'hB5;
                    16'hE5D1: data_out = 8'hB6;
                    16'hE5D2: data_out = 8'hB7;
                    16'hE5D3: data_out = 8'hB8;
                    16'hE5D4: data_out = 8'hB9;
                    16'hE5D5: data_out = 8'hBA;
                    16'hE5D6: data_out = 8'hBB;
                    16'hE5D7: data_out = 8'hBC;
                    16'hE5D8: data_out = 8'hBD;
                    16'hE5D9: data_out = 8'hBE;
                    16'hE5DA: data_out = 8'hBF;
                    16'hE5DB: data_out = 8'hC0;
                    16'hE5DC: data_out = 8'hC1;
                    16'hE5DD: data_out = 8'hC2;
                    16'hE5DE: data_out = 8'hC3;
                    16'hE5DF: data_out = 8'hC4;
                    16'hE5E0: data_out = 8'hC5;
                    16'hE5E1: data_out = 8'hC6;
                    16'hE5E2: data_out = 8'hC7;
                    16'hE5E3: data_out = 8'hC8;
                    16'hE5E4: data_out = 8'hC9;
                    16'hE5E5: data_out = 8'hCA;
                    16'hE5E6: data_out = 8'hCB;
                    16'hE5E7: data_out = 8'hCC;
                    16'hE5E8: data_out = 8'hCD;
                    16'hE5E9: data_out = 8'hCE;
                    16'hE5EA: data_out = 8'hCF;
                    16'hE5EB: data_out = 8'hD0;
                    16'hE5EC: data_out = 8'hD1;
                    16'hE5ED: data_out = 8'hD2;
                    16'hE5EE: data_out = 8'hD3;
                    16'hE5EF: data_out = 8'hD4;
                    16'hE5F0: data_out = 8'hD5;
                    16'hE5F1: data_out = 8'hD6;
                    16'hE5F2: data_out = 8'hD7;
                    16'hE5F3: data_out = 8'hD8;
                    16'hE5F4: data_out = 8'hD9;
                    16'hE5F5: data_out = 8'hDA;
                    16'hE5F6: data_out = 8'hDB;
                    16'hE5F7: data_out = 8'hDC;
                    16'hE5F8: data_out = 8'hDD;
                    16'hE5F9: data_out = 8'hDE;
                    16'hE5FA: data_out = 8'hDF;
                    16'hE5FB: data_out = 8'hE0;
                    16'hE5FC: data_out = 8'hE1;
                    16'hE5FD: data_out = 8'hE2;
                    16'hE5FE: data_out = 8'hE3;
                    16'hE5FF: data_out = 8'hE4;
                    16'hE600: data_out = 8'hE6;
                    16'hE601: data_out = 8'hE5;
                    16'hE602: data_out = 8'hE4;
                    16'hE603: data_out = 8'hE3;
                    16'hE604: data_out = 8'hE2;
                    16'hE605: data_out = 8'hE1;
                    16'hE606: data_out = 8'hE0;
                    16'hE607: data_out = 8'hDF;
                    16'hE608: data_out = 8'hDE;
                    16'hE609: data_out = 8'hDD;
                    16'hE60A: data_out = 8'hDC;
                    16'hE60B: data_out = 8'hDB;
                    16'hE60C: data_out = 8'hDA;
                    16'hE60D: data_out = 8'hD9;
                    16'hE60E: data_out = 8'hD8;
                    16'hE60F: data_out = 8'hD7;
                    16'hE610: data_out = 8'hD6;
                    16'hE611: data_out = 8'hD5;
                    16'hE612: data_out = 8'hD4;
                    16'hE613: data_out = 8'hD3;
                    16'hE614: data_out = 8'hD2;
                    16'hE615: data_out = 8'hD1;
                    16'hE616: data_out = 8'hD0;
                    16'hE617: data_out = 8'hCF;
                    16'hE618: data_out = 8'hCE;
                    16'hE619: data_out = 8'hCD;
                    16'hE61A: data_out = 8'hCC;
                    16'hE61B: data_out = 8'hCB;
                    16'hE61C: data_out = 8'hCA;
                    16'hE61D: data_out = 8'hC9;
                    16'hE61E: data_out = 8'hC8;
                    16'hE61F: data_out = 8'hC7;
                    16'hE620: data_out = 8'hC6;
                    16'hE621: data_out = 8'hC5;
                    16'hE622: data_out = 8'hC4;
                    16'hE623: data_out = 8'hC3;
                    16'hE624: data_out = 8'hC2;
                    16'hE625: data_out = 8'hC1;
                    16'hE626: data_out = 8'hC0;
                    16'hE627: data_out = 8'hBF;
                    16'hE628: data_out = 8'hBE;
                    16'hE629: data_out = 8'hBD;
                    16'hE62A: data_out = 8'hBC;
                    16'hE62B: data_out = 8'hBB;
                    16'hE62C: data_out = 8'hBA;
                    16'hE62D: data_out = 8'hB9;
                    16'hE62E: data_out = 8'hB8;
                    16'hE62F: data_out = 8'hB7;
                    16'hE630: data_out = 8'hB6;
                    16'hE631: data_out = 8'hB5;
                    16'hE632: data_out = 8'hB4;
                    16'hE633: data_out = 8'hB3;
                    16'hE634: data_out = 8'hB2;
                    16'hE635: data_out = 8'hB1;
                    16'hE636: data_out = 8'hB0;
                    16'hE637: data_out = 8'hAF;
                    16'hE638: data_out = 8'hAE;
                    16'hE639: data_out = 8'hAD;
                    16'hE63A: data_out = 8'hAC;
                    16'hE63B: data_out = 8'hAB;
                    16'hE63C: data_out = 8'hAA;
                    16'hE63D: data_out = 8'hA9;
                    16'hE63E: data_out = 8'hA8;
                    16'hE63F: data_out = 8'hA7;
                    16'hE640: data_out = 8'hA6;
                    16'hE641: data_out = 8'hA5;
                    16'hE642: data_out = 8'hA4;
                    16'hE643: data_out = 8'hA3;
                    16'hE644: data_out = 8'hA2;
                    16'hE645: data_out = 8'hA1;
                    16'hE646: data_out = 8'hA0;
                    16'hE647: data_out = 8'h9F;
                    16'hE648: data_out = 8'h9E;
                    16'hE649: data_out = 8'h9D;
                    16'hE64A: data_out = 8'h9C;
                    16'hE64B: data_out = 8'h9B;
                    16'hE64C: data_out = 8'h9A;
                    16'hE64D: data_out = 8'h99;
                    16'hE64E: data_out = 8'h98;
                    16'hE64F: data_out = 8'h97;
                    16'hE650: data_out = 8'h96;
                    16'hE651: data_out = 8'h95;
                    16'hE652: data_out = 8'h94;
                    16'hE653: data_out = 8'h93;
                    16'hE654: data_out = 8'h92;
                    16'hE655: data_out = 8'h91;
                    16'hE656: data_out = 8'h90;
                    16'hE657: data_out = 8'h8F;
                    16'hE658: data_out = 8'h8E;
                    16'hE659: data_out = 8'h8D;
                    16'hE65A: data_out = 8'h8C;
                    16'hE65B: data_out = 8'h8B;
                    16'hE65C: data_out = 8'h8A;
                    16'hE65D: data_out = 8'h89;
                    16'hE65E: data_out = 8'h88;
                    16'hE65F: data_out = 8'h87;
                    16'hE660: data_out = 8'h86;
                    16'hE661: data_out = 8'h85;
                    16'hE662: data_out = 8'h84;
                    16'hE663: data_out = 8'h83;
                    16'hE664: data_out = 8'h82;
                    16'hE665: data_out = 8'h81;
                    16'hE666: data_out = 8'h0;
                    16'hE667: data_out = 8'h1;
                    16'hE668: data_out = 8'h2;
                    16'hE669: data_out = 8'h3;
                    16'hE66A: data_out = 8'h4;
                    16'hE66B: data_out = 8'h5;
                    16'hE66C: data_out = 8'h6;
                    16'hE66D: data_out = 8'h7;
                    16'hE66E: data_out = 8'h8;
                    16'hE66F: data_out = 8'h9;
                    16'hE670: data_out = 8'hA;
                    16'hE671: data_out = 8'hB;
                    16'hE672: data_out = 8'hC;
                    16'hE673: data_out = 8'hD;
                    16'hE674: data_out = 8'hE;
                    16'hE675: data_out = 8'hF;
                    16'hE676: data_out = 8'h10;
                    16'hE677: data_out = 8'h11;
                    16'hE678: data_out = 8'h12;
                    16'hE679: data_out = 8'h13;
                    16'hE67A: data_out = 8'h14;
                    16'hE67B: data_out = 8'h15;
                    16'hE67C: data_out = 8'h16;
                    16'hE67D: data_out = 8'h17;
                    16'hE67E: data_out = 8'h18;
                    16'hE67F: data_out = 8'h19;
                    16'hE680: data_out = 8'hE6;
                    16'hE681: data_out = 8'hE7;
                    16'hE682: data_out = 8'hE8;
                    16'hE683: data_out = 8'hE9;
                    16'hE684: data_out = 8'hEA;
                    16'hE685: data_out = 8'hEB;
                    16'hE686: data_out = 8'hEC;
                    16'hE687: data_out = 8'hED;
                    16'hE688: data_out = 8'hEE;
                    16'hE689: data_out = 8'hEF;
                    16'hE68A: data_out = 8'hF0;
                    16'hE68B: data_out = 8'hF1;
                    16'hE68C: data_out = 8'hF2;
                    16'hE68D: data_out = 8'hF3;
                    16'hE68E: data_out = 8'hF4;
                    16'hE68F: data_out = 8'hF5;
                    16'hE690: data_out = 8'hF6;
                    16'hE691: data_out = 8'hF7;
                    16'hE692: data_out = 8'hF8;
                    16'hE693: data_out = 8'hF9;
                    16'hE694: data_out = 8'hFA;
                    16'hE695: data_out = 8'hFB;
                    16'hE696: data_out = 8'hFC;
                    16'hE697: data_out = 8'hFD;
                    16'hE698: data_out = 8'hFE;
                    16'hE699: data_out = 8'hFF;
                    16'hE69A: data_out = 8'h80;
                    16'hE69B: data_out = 8'h81;
                    16'hE69C: data_out = 8'h82;
                    16'hE69D: data_out = 8'h83;
                    16'hE69E: data_out = 8'h84;
                    16'hE69F: data_out = 8'h85;
                    16'hE6A0: data_out = 8'h86;
                    16'hE6A1: data_out = 8'h87;
                    16'hE6A2: data_out = 8'h88;
                    16'hE6A3: data_out = 8'h89;
                    16'hE6A4: data_out = 8'h8A;
                    16'hE6A5: data_out = 8'h8B;
                    16'hE6A6: data_out = 8'h8C;
                    16'hE6A7: data_out = 8'h8D;
                    16'hE6A8: data_out = 8'h8E;
                    16'hE6A9: data_out = 8'h8F;
                    16'hE6AA: data_out = 8'h90;
                    16'hE6AB: data_out = 8'h91;
                    16'hE6AC: data_out = 8'h92;
                    16'hE6AD: data_out = 8'h93;
                    16'hE6AE: data_out = 8'h94;
                    16'hE6AF: data_out = 8'h95;
                    16'hE6B0: data_out = 8'h96;
                    16'hE6B1: data_out = 8'h97;
                    16'hE6B2: data_out = 8'h98;
                    16'hE6B3: data_out = 8'h99;
                    16'hE6B4: data_out = 8'h9A;
                    16'hE6B5: data_out = 8'h9B;
                    16'hE6B6: data_out = 8'h9C;
                    16'hE6B7: data_out = 8'h9D;
                    16'hE6B8: data_out = 8'h9E;
                    16'hE6B9: data_out = 8'h9F;
                    16'hE6BA: data_out = 8'hA0;
                    16'hE6BB: data_out = 8'hA1;
                    16'hE6BC: data_out = 8'hA2;
                    16'hE6BD: data_out = 8'hA3;
                    16'hE6BE: data_out = 8'hA4;
                    16'hE6BF: data_out = 8'hA5;
                    16'hE6C0: data_out = 8'hA6;
                    16'hE6C1: data_out = 8'hA7;
                    16'hE6C2: data_out = 8'hA8;
                    16'hE6C3: data_out = 8'hA9;
                    16'hE6C4: data_out = 8'hAA;
                    16'hE6C5: data_out = 8'hAB;
                    16'hE6C6: data_out = 8'hAC;
                    16'hE6C7: data_out = 8'hAD;
                    16'hE6C8: data_out = 8'hAE;
                    16'hE6C9: data_out = 8'hAF;
                    16'hE6CA: data_out = 8'hB0;
                    16'hE6CB: data_out = 8'hB1;
                    16'hE6CC: data_out = 8'hB2;
                    16'hE6CD: data_out = 8'hB3;
                    16'hE6CE: data_out = 8'hB4;
                    16'hE6CF: data_out = 8'hB5;
                    16'hE6D0: data_out = 8'hB6;
                    16'hE6D1: data_out = 8'hB7;
                    16'hE6D2: data_out = 8'hB8;
                    16'hE6D3: data_out = 8'hB9;
                    16'hE6D4: data_out = 8'hBA;
                    16'hE6D5: data_out = 8'hBB;
                    16'hE6D6: data_out = 8'hBC;
                    16'hE6D7: data_out = 8'hBD;
                    16'hE6D8: data_out = 8'hBE;
                    16'hE6D9: data_out = 8'hBF;
                    16'hE6DA: data_out = 8'hC0;
                    16'hE6DB: data_out = 8'hC1;
                    16'hE6DC: data_out = 8'hC2;
                    16'hE6DD: data_out = 8'hC3;
                    16'hE6DE: data_out = 8'hC4;
                    16'hE6DF: data_out = 8'hC5;
                    16'hE6E0: data_out = 8'hC6;
                    16'hE6E1: data_out = 8'hC7;
                    16'hE6E2: data_out = 8'hC8;
                    16'hE6E3: data_out = 8'hC9;
                    16'hE6E4: data_out = 8'hCA;
                    16'hE6E5: data_out = 8'hCB;
                    16'hE6E6: data_out = 8'hCC;
                    16'hE6E7: data_out = 8'hCD;
                    16'hE6E8: data_out = 8'hCE;
                    16'hE6E9: data_out = 8'hCF;
                    16'hE6EA: data_out = 8'hD0;
                    16'hE6EB: data_out = 8'hD1;
                    16'hE6EC: data_out = 8'hD2;
                    16'hE6ED: data_out = 8'hD3;
                    16'hE6EE: data_out = 8'hD4;
                    16'hE6EF: data_out = 8'hD5;
                    16'hE6F0: data_out = 8'hD6;
                    16'hE6F1: data_out = 8'hD7;
                    16'hE6F2: data_out = 8'hD8;
                    16'hE6F3: data_out = 8'hD9;
                    16'hE6F4: data_out = 8'hDA;
                    16'hE6F5: data_out = 8'hDB;
                    16'hE6F6: data_out = 8'hDC;
                    16'hE6F7: data_out = 8'hDD;
                    16'hE6F8: data_out = 8'hDE;
                    16'hE6F9: data_out = 8'hDF;
                    16'hE6FA: data_out = 8'hE0;
                    16'hE6FB: data_out = 8'hE1;
                    16'hE6FC: data_out = 8'hE2;
                    16'hE6FD: data_out = 8'hE3;
                    16'hE6FE: data_out = 8'hE4;
                    16'hE6FF: data_out = 8'hE5;
                    16'hE700: data_out = 8'hE7;
                    16'hE701: data_out = 8'hE6;
                    16'hE702: data_out = 8'hE5;
                    16'hE703: data_out = 8'hE4;
                    16'hE704: data_out = 8'hE3;
                    16'hE705: data_out = 8'hE2;
                    16'hE706: data_out = 8'hE1;
                    16'hE707: data_out = 8'hE0;
                    16'hE708: data_out = 8'hDF;
                    16'hE709: data_out = 8'hDE;
                    16'hE70A: data_out = 8'hDD;
                    16'hE70B: data_out = 8'hDC;
                    16'hE70C: data_out = 8'hDB;
                    16'hE70D: data_out = 8'hDA;
                    16'hE70E: data_out = 8'hD9;
                    16'hE70F: data_out = 8'hD8;
                    16'hE710: data_out = 8'hD7;
                    16'hE711: data_out = 8'hD6;
                    16'hE712: data_out = 8'hD5;
                    16'hE713: data_out = 8'hD4;
                    16'hE714: data_out = 8'hD3;
                    16'hE715: data_out = 8'hD2;
                    16'hE716: data_out = 8'hD1;
                    16'hE717: data_out = 8'hD0;
                    16'hE718: data_out = 8'hCF;
                    16'hE719: data_out = 8'hCE;
                    16'hE71A: data_out = 8'hCD;
                    16'hE71B: data_out = 8'hCC;
                    16'hE71C: data_out = 8'hCB;
                    16'hE71D: data_out = 8'hCA;
                    16'hE71E: data_out = 8'hC9;
                    16'hE71F: data_out = 8'hC8;
                    16'hE720: data_out = 8'hC7;
                    16'hE721: data_out = 8'hC6;
                    16'hE722: data_out = 8'hC5;
                    16'hE723: data_out = 8'hC4;
                    16'hE724: data_out = 8'hC3;
                    16'hE725: data_out = 8'hC2;
                    16'hE726: data_out = 8'hC1;
                    16'hE727: data_out = 8'hC0;
                    16'hE728: data_out = 8'hBF;
                    16'hE729: data_out = 8'hBE;
                    16'hE72A: data_out = 8'hBD;
                    16'hE72B: data_out = 8'hBC;
                    16'hE72C: data_out = 8'hBB;
                    16'hE72D: data_out = 8'hBA;
                    16'hE72E: data_out = 8'hB9;
                    16'hE72F: data_out = 8'hB8;
                    16'hE730: data_out = 8'hB7;
                    16'hE731: data_out = 8'hB6;
                    16'hE732: data_out = 8'hB5;
                    16'hE733: data_out = 8'hB4;
                    16'hE734: data_out = 8'hB3;
                    16'hE735: data_out = 8'hB2;
                    16'hE736: data_out = 8'hB1;
                    16'hE737: data_out = 8'hB0;
                    16'hE738: data_out = 8'hAF;
                    16'hE739: data_out = 8'hAE;
                    16'hE73A: data_out = 8'hAD;
                    16'hE73B: data_out = 8'hAC;
                    16'hE73C: data_out = 8'hAB;
                    16'hE73D: data_out = 8'hAA;
                    16'hE73E: data_out = 8'hA9;
                    16'hE73F: data_out = 8'hA8;
                    16'hE740: data_out = 8'hA7;
                    16'hE741: data_out = 8'hA6;
                    16'hE742: data_out = 8'hA5;
                    16'hE743: data_out = 8'hA4;
                    16'hE744: data_out = 8'hA3;
                    16'hE745: data_out = 8'hA2;
                    16'hE746: data_out = 8'hA1;
                    16'hE747: data_out = 8'hA0;
                    16'hE748: data_out = 8'h9F;
                    16'hE749: data_out = 8'h9E;
                    16'hE74A: data_out = 8'h9D;
                    16'hE74B: data_out = 8'h9C;
                    16'hE74C: data_out = 8'h9B;
                    16'hE74D: data_out = 8'h9A;
                    16'hE74E: data_out = 8'h99;
                    16'hE74F: data_out = 8'h98;
                    16'hE750: data_out = 8'h97;
                    16'hE751: data_out = 8'h96;
                    16'hE752: data_out = 8'h95;
                    16'hE753: data_out = 8'h94;
                    16'hE754: data_out = 8'h93;
                    16'hE755: data_out = 8'h92;
                    16'hE756: data_out = 8'h91;
                    16'hE757: data_out = 8'h90;
                    16'hE758: data_out = 8'h8F;
                    16'hE759: data_out = 8'h8E;
                    16'hE75A: data_out = 8'h8D;
                    16'hE75B: data_out = 8'h8C;
                    16'hE75C: data_out = 8'h8B;
                    16'hE75D: data_out = 8'h8A;
                    16'hE75E: data_out = 8'h89;
                    16'hE75F: data_out = 8'h88;
                    16'hE760: data_out = 8'h87;
                    16'hE761: data_out = 8'h86;
                    16'hE762: data_out = 8'h85;
                    16'hE763: data_out = 8'h84;
                    16'hE764: data_out = 8'h83;
                    16'hE765: data_out = 8'h82;
                    16'hE766: data_out = 8'h81;
                    16'hE767: data_out = 8'h0;
                    16'hE768: data_out = 8'h1;
                    16'hE769: data_out = 8'h2;
                    16'hE76A: data_out = 8'h3;
                    16'hE76B: data_out = 8'h4;
                    16'hE76C: data_out = 8'h5;
                    16'hE76D: data_out = 8'h6;
                    16'hE76E: data_out = 8'h7;
                    16'hE76F: data_out = 8'h8;
                    16'hE770: data_out = 8'h9;
                    16'hE771: data_out = 8'hA;
                    16'hE772: data_out = 8'hB;
                    16'hE773: data_out = 8'hC;
                    16'hE774: data_out = 8'hD;
                    16'hE775: data_out = 8'hE;
                    16'hE776: data_out = 8'hF;
                    16'hE777: data_out = 8'h10;
                    16'hE778: data_out = 8'h11;
                    16'hE779: data_out = 8'h12;
                    16'hE77A: data_out = 8'h13;
                    16'hE77B: data_out = 8'h14;
                    16'hE77C: data_out = 8'h15;
                    16'hE77D: data_out = 8'h16;
                    16'hE77E: data_out = 8'h17;
                    16'hE77F: data_out = 8'h18;
                    16'hE780: data_out = 8'hE7;
                    16'hE781: data_out = 8'hE8;
                    16'hE782: data_out = 8'hE9;
                    16'hE783: data_out = 8'hEA;
                    16'hE784: data_out = 8'hEB;
                    16'hE785: data_out = 8'hEC;
                    16'hE786: data_out = 8'hED;
                    16'hE787: data_out = 8'hEE;
                    16'hE788: data_out = 8'hEF;
                    16'hE789: data_out = 8'hF0;
                    16'hE78A: data_out = 8'hF1;
                    16'hE78B: data_out = 8'hF2;
                    16'hE78C: data_out = 8'hF3;
                    16'hE78D: data_out = 8'hF4;
                    16'hE78E: data_out = 8'hF5;
                    16'hE78F: data_out = 8'hF6;
                    16'hE790: data_out = 8'hF7;
                    16'hE791: data_out = 8'hF8;
                    16'hE792: data_out = 8'hF9;
                    16'hE793: data_out = 8'hFA;
                    16'hE794: data_out = 8'hFB;
                    16'hE795: data_out = 8'hFC;
                    16'hE796: data_out = 8'hFD;
                    16'hE797: data_out = 8'hFE;
                    16'hE798: data_out = 8'hFF;
                    16'hE799: data_out = 8'h80;
                    16'hE79A: data_out = 8'h81;
                    16'hE79B: data_out = 8'h82;
                    16'hE79C: data_out = 8'h83;
                    16'hE79D: data_out = 8'h84;
                    16'hE79E: data_out = 8'h85;
                    16'hE79F: data_out = 8'h86;
                    16'hE7A0: data_out = 8'h87;
                    16'hE7A1: data_out = 8'h88;
                    16'hE7A2: data_out = 8'h89;
                    16'hE7A3: data_out = 8'h8A;
                    16'hE7A4: data_out = 8'h8B;
                    16'hE7A5: data_out = 8'h8C;
                    16'hE7A6: data_out = 8'h8D;
                    16'hE7A7: data_out = 8'h8E;
                    16'hE7A8: data_out = 8'h8F;
                    16'hE7A9: data_out = 8'h90;
                    16'hE7AA: data_out = 8'h91;
                    16'hE7AB: data_out = 8'h92;
                    16'hE7AC: data_out = 8'h93;
                    16'hE7AD: data_out = 8'h94;
                    16'hE7AE: data_out = 8'h95;
                    16'hE7AF: data_out = 8'h96;
                    16'hE7B0: data_out = 8'h97;
                    16'hE7B1: data_out = 8'h98;
                    16'hE7B2: data_out = 8'h99;
                    16'hE7B3: data_out = 8'h9A;
                    16'hE7B4: data_out = 8'h9B;
                    16'hE7B5: data_out = 8'h9C;
                    16'hE7B6: data_out = 8'h9D;
                    16'hE7B7: data_out = 8'h9E;
                    16'hE7B8: data_out = 8'h9F;
                    16'hE7B9: data_out = 8'hA0;
                    16'hE7BA: data_out = 8'hA1;
                    16'hE7BB: data_out = 8'hA2;
                    16'hE7BC: data_out = 8'hA3;
                    16'hE7BD: data_out = 8'hA4;
                    16'hE7BE: data_out = 8'hA5;
                    16'hE7BF: data_out = 8'hA6;
                    16'hE7C0: data_out = 8'hA7;
                    16'hE7C1: data_out = 8'hA8;
                    16'hE7C2: data_out = 8'hA9;
                    16'hE7C3: data_out = 8'hAA;
                    16'hE7C4: data_out = 8'hAB;
                    16'hE7C5: data_out = 8'hAC;
                    16'hE7C6: data_out = 8'hAD;
                    16'hE7C7: data_out = 8'hAE;
                    16'hE7C8: data_out = 8'hAF;
                    16'hE7C9: data_out = 8'hB0;
                    16'hE7CA: data_out = 8'hB1;
                    16'hE7CB: data_out = 8'hB2;
                    16'hE7CC: data_out = 8'hB3;
                    16'hE7CD: data_out = 8'hB4;
                    16'hE7CE: data_out = 8'hB5;
                    16'hE7CF: data_out = 8'hB6;
                    16'hE7D0: data_out = 8'hB7;
                    16'hE7D1: data_out = 8'hB8;
                    16'hE7D2: data_out = 8'hB9;
                    16'hE7D3: data_out = 8'hBA;
                    16'hE7D4: data_out = 8'hBB;
                    16'hE7D5: data_out = 8'hBC;
                    16'hE7D6: data_out = 8'hBD;
                    16'hE7D7: data_out = 8'hBE;
                    16'hE7D8: data_out = 8'hBF;
                    16'hE7D9: data_out = 8'hC0;
                    16'hE7DA: data_out = 8'hC1;
                    16'hE7DB: data_out = 8'hC2;
                    16'hE7DC: data_out = 8'hC3;
                    16'hE7DD: data_out = 8'hC4;
                    16'hE7DE: data_out = 8'hC5;
                    16'hE7DF: data_out = 8'hC6;
                    16'hE7E0: data_out = 8'hC7;
                    16'hE7E1: data_out = 8'hC8;
                    16'hE7E2: data_out = 8'hC9;
                    16'hE7E3: data_out = 8'hCA;
                    16'hE7E4: data_out = 8'hCB;
                    16'hE7E5: data_out = 8'hCC;
                    16'hE7E6: data_out = 8'hCD;
                    16'hE7E7: data_out = 8'hCE;
                    16'hE7E8: data_out = 8'hCF;
                    16'hE7E9: data_out = 8'hD0;
                    16'hE7EA: data_out = 8'hD1;
                    16'hE7EB: data_out = 8'hD2;
                    16'hE7EC: data_out = 8'hD3;
                    16'hE7ED: data_out = 8'hD4;
                    16'hE7EE: data_out = 8'hD5;
                    16'hE7EF: data_out = 8'hD6;
                    16'hE7F0: data_out = 8'hD7;
                    16'hE7F1: data_out = 8'hD8;
                    16'hE7F2: data_out = 8'hD9;
                    16'hE7F3: data_out = 8'hDA;
                    16'hE7F4: data_out = 8'hDB;
                    16'hE7F5: data_out = 8'hDC;
                    16'hE7F6: data_out = 8'hDD;
                    16'hE7F7: data_out = 8'hDE;
                    16'hE7F8: data_out = 8'hDF;
                    16'hE7F9: data_out = 8'hE0;
                    16'hE7FA: data_out = 8'hE1;
                    16'hE7FB: data_out = 8'hE2;
                    16'hE7FC: data_out = 8'hE3;
                    16'hE7FD: data_out = 8'hE4;
                    16'hE7FE: data_out = 8'hE5;
                    16'hE7FF: data_out = 8'hE6;
                    16'hE800: data_out = 8'hE8;
                    16'hE801: data_out = 8'hE7;
                    16'hE802: data_out = 8'hE6;
                    16'hE803: data_out = 8'hE5;
                    16'hE804: data_out = 8'hE4;
                    16'hE805: data_out = 8'hE3;
                    16'hE806: data_out = 8'hE2;
                    16'hE807: data_out = 8'hE1;
                    16'hE808: data_out = 8'hE0;
                    16'hE809: data_out = 8'hDF;
                    16'hE80A: data_out = 8'hDE;
                    16'hE80B: data_out = 8'hDD;
                    16'hE80C: data_out = 8'hDC;
                    16'hE80D: data_out = 8'hDB;
                    16'hE80E: data_out = 8'hDA;
                    16'hE80F: data_out = 8'hD9;
                    16'hE810: data_out = 8'hD8;
                    16'hE811: data_out = 8'hD7;
                    16'hE812: data_out = 8'hD6;
                    16'hE813: data_out = 8'hD5;
                    16'hE814: data_out = 8'hD4;
                    16'hE815: data_out = 8'hD3;
                    16'hE816: data_out = 8'hD2;
                    16'hE817: data_out = 8'hD1;
                    16'hE818: data_out = 8'hD0;
                    16'hE819: data_out = 8'hCF;
                    16'hE81A: data_out = 8'hCE;
                    16'hE81B: data_out = 8'hCD;
                    16'hE81C: data_out = 8'hCC;
                    16'hE81D: data_out = 8'hCB;
                    16'hE81E: data_out = 8'hCA;
                    16'hE81F: data_out = 8'hC9;
                    16'hE820: data_out = 8'hC8;
                    16'hE821: data_out = 8'hC7;
                    16'hE822: data_out = 8'hC6;
                    16'hE823: data_out = 8'hC5;
                    16'hE824: data_out = 8'hC4;
                    16'hE825: data_out = 8'hC3;
                    16'hE826: data_out = 8'hC2;
                    16'hE827: data_out = 8'hC1;
                    16'hE828: data_out = 8'hC0;
                    16'hE829: data_out = 8'hBF;
                    16'hE82A: data_out = 8'hBE;
                    16'hE82B: data_out = 8'hBD;
                    16'hE82C: data_out = 8'hBC;
                    16'hE82D: data_out = 8'hBB;
                    16'hE82E: data_out = 8'hBA;
                    16'hE82F: data_out = 8'hB9;
                    16'hE830: data_out = 8'hB8;
                    16'hE831: data_out = 8'hB7;
                    16'hE832: data_out = 8'hB6;
                    16'hE833: data_out = 8'hB5;
                    16'hE834: data_out = 8'hB4;
                    16'hE835: data_out = 8'hB3;
                    16'hE836: data_out = 8'hB2;
                    16'hE837: data_out = 8'hB1;
                    16'hE838: data_out = 8'hB0;
                    16'hE839: data_out = 8'hAF;
                    16'hE83A: data_out = 8'hAE;
                    16'hE83B: data_out = 8'hAD;
                    16'hE83C: data_out = 8'hAC;
                    16'hE83D: data_out = 8'hAB;
                    16'hE83E: data_out = 8'hAA;
                    16'hE83F: data_out = 8'hA9;
                    16'hE840: data_out = 8'hA8;
                    16'hE841: data_out = 8'hA7;
                    16'hE842: data_out = 8'hA6;
                    16'hE843: data_out = 8'hA5;
                    16'hE844: data_out = 8'hA4;
                    16'hE845: data_out = 8'hA3;
                    16'hE846: data_out = 8'hA2;
                    16'hE847: data_out = 8'hA1;
                    16'hE848: data_out = 8'hA0;
                    16'hE849: data_out = 8'h9F;
                    16'hE84A: data_out = 8'h9E;
                    16'hE84B: data_out = 8'h9D;
                    16'hE84C: data_out = 8'h9C;
                    16'hE84D: data_out = 8'h9B;
                    16'hE84E: data_out = 8'h9A;
                    16'hE84F: data_out = 8'h99;
                    16'hE850: data_out = 8'h98;
                    16'hE851: data_out = 8'h97;
                    16'hE852: data_out = 8'h96;
                    16'hE853: data_out = 8'h95;
                    16'hE854: data_out = 8'h94;
                    16'hE855: data_out = 8'h93;
                    16'hE856: data_out = 8'h92;
                    16'hE857: data_out = 8'h91;
                    16'hE858: data_out = 8'h90;
                    16'hE859: data_out = 8'h8F;
                    16'hE85A: data_out = 8'h8E;
                    16'hE85B: data_out = 8'h8D;
                    16'hE85C: data_out = 8'h8C;
                    16'hE85D: data_out = 8'h8B;
                    16'hE85E: data_out = 8'h8A;
                    16'hE85F: data_out = 8'h89;
                    16'hE860: data_out = 8'h88;
                    16'hE861: data_out = 8'h87;
                    16'hE862: data_out = 8'h86;
                    16'hE863: data_out = 8'h85;
                    16'hE864: data_out = 8'h84;
                    16'hE865: data_out = 8'h83;
                    16'hE866: data_out = 8'h82;
                    16'hE867: data_out = 8'h81;
                    16'hE868: data_out = 8'h0;
                    16'hE869: data_out = 8'h1;
                    16'hE86A: data_out = 8'h2;
                    16'hE86B: data_out = 8'h3;
                    16'hE86C: data_out = 8'h4;
                    16'hE86D: data_out = 8'h5;
                    16'hE86E: data_out = 8'h6;
                    16'hE86F: data_out = 8'h7;
                    16'hE870: data_out = 8'h8;
                    16'hE871: data_out = 8'h9;
                    16'hE872: data_out = 8'hA;
                    16'hE873: data_out = 8'hB;
                    16'hE874: data_out = 8'hC;
                    16'hE875: data_out = 8'hD;
                    16'hE876: data_out = 8'hE;
                    16'hE877: data_out = 8'hF;
                    16'hE878: data_out = 8'h10;
                    16'hE879: data_out = 8'h11;
                    16'hE87A: data_out = 8'h12;
                    16'hE87B: data_out = 8'h13;
                    16'hE87C: data_out = 8'h14;
                    16'hE87D: data_out = 8'h15;
                    16'hE87E: data_out = 8'h16;
                    16'hE87F: data_out = 8'h17;
                    16'hE880: data_out = 8'hE8;
                    16'hE881: data_out = 8'hE9;
                    16'hE882: data_out = 8'hEA;
                    16'hE883: data_out = 8'hEB;
                    16'hE884: data_out = 8'hEC;
                    16'hE885: data_out = 8'hED;
                    16'hE886: data_out = 8'hEE;
                    16'hE887: data_out = 8'hEF;
                    16'hE888: data_out = 8'hF0;
                    16'hE889: data_out = 8'hF1;
                    16'hE88A: data_out = 8'hF2;
                    16'hE88B: data_out = 8'hF3;
                    16'hE88C: data_out = 8'hF4;
                    16'hE88D: data_out = 8'hF5;
                    16'hE88E: data_out = 8'hF6;
                    16'hE88F: data_out = 8'hF7;
                    16'hE890: data_out = 8'hF8;
                    16'hE891: data_out = 8'hF9;
                    16'hE892: data_out = 8'hFA;
                    16'hE893: data_out = 8'hFB;
                    16'hE894: data_out = 8'hFC;
                    16'hE895: data_out = 8'hFD;
                    16'hE896: data_out = 8'hFE;
                    16'hE897: data_out = 8'hFF;
                    16'hE898: data_out = 8'h80;
                    16'hE899: data_out = 8'h81;
                    16'hE89A: data_out = 8'h82;
                    16'hE89B: data_out = 8'h83;
                    16'hE89C: data_out = 8'h84;
                    16'hE89D: data_out = 8'h85;
                    16'hE89E: data_out = 8'h86;
                    16'hE89F: data_out = 8'h87;
                    16'hE8A0: data_out = 8'h88;
                    16'hE8A1: data_out = 8'h89;
                    16'hE8A2: data_out = 8'h8A;
                    16'hE8A3: data_out = 8'h8B;
                    16'hE8A4: data_out = 8'h8C;
                    16'hE8A5: data_out = 8'h8D;
                    16'hE8A6: data_out = 8'h8E;
                    16'hE8A7: data_out = 8'h8F;
                    16'hE8A8: data_out = 8'h90;
                    16'hE8A9: data_out = 8'h91;
                    16'hE8AA: data_out = 8'h92;
                    16'hE8AB: data_out = 8'h93;
                    16'hE8AC: data_out = 8'h94;
                    16'hE8AD: data_out = 8'h95;
                    16'hE8AE: data_out = 8'h96;
                    16'hE8AF: data_out = 8'h97;
                    16'hE8B0: data_out = 8'h98;
                    16'hE8B1: data_out = 8'h99;
                    16'hE8B2: data_out = 8'h9A;
                    16'hE8B3: data_out = 8'h9B;
                    16'hE8B4: data_out = 8'h9C;
                    16'hE8B5: data_out = 8'h9D;
                    16'hE8B6: data_out = 8'h9E;
                    16'hE8B7: data_out = 8'h9F;
                    16'hE8B8: data_out = 8'hA0;
                    16'hE8B9: data_out = 8'hA1;
                    16'hE8BA: data_out = 8'hA2;
                    16'hE8BB: data_out = 8'hA3;
                    16'hE8BC: data_out = 8'hA4;
                    16'hE8BD: data_out = 8'hA5;
                    16'hE8BE: data_out = 8'hA6;
                    16'hE8BF: data_out = 8'hA7;
                    16'hE8C0: data_out = 8'hA8;
                    16'hE8C1: data_out = 8'hA9;
                    16'hE8C2: data_out = 8'hAA;
                    16'hE8C3: data_out = 8'hAB;
                    16'hE8C4: data_out = 8'hAC;
                    16'hE8C5: data_out = 8'hAD;
                    16'hE8C6: data_out = 8'hAE;
                    16'hE8C7: data_out = 8'hAF;
                    16'hE8C8: data_out = 8'hB0;
                    16'hE8C9: data_out = 8'hB1;
                    16'hE8CA: data_out = 8'hB2;
                    16'hE8CB: data_out = 8'hB3;
                    16'hE8CC: data_out = 8'hB4;
                    16'hE8CD: data_out = 8'hB5;
                    16'hE8CE: data_out = 8'hB6;
                    16'hE8CF: data_out = 8'hB7;
                    16'hE8D0: data_out = 8'hB8;
                    16'hE8D1: data_out = 8'hB9;
                    16'hE8D2: data_out = 8'hBA;
                    16'hE8D3: data_out = 8'hBB;
                    16'hE8D4: data_out = 8'hBC;
                    16'hE8D5: data_out = 8'hBD;
                    16'hE8D6: data_out = 8'hBE;
                    16'hE8D7: data_out = 8'hBF;
                    16'hE8D8: data_out = 8'hC0;
                    16'hE8D9: data_out = 8'hC1;
                    16'hE8DA: data_out = 8'hC2;
                    16'hE8DB: data_out = 8'hC3;
                    16'hE8DC: data_out = 8'hC4;
                    16'hE8DD: data_out = 8'hC5;
                    16'hE8DE: data_out = 8'hC6;
                    16'hE8DF: data_out = 8'hC7;
                    16'hE8E0: data_out = 8'hC8;
                    16'hE8E1: data_out = 8'hC9;
                    16'hE8E2: data_out = 8'hCA;
                    16'hE8E3: data_out = 8'hCB;
                    16'hE8E4: data_out = 8'hCC;
                    16'hE8E5: data_out = 8'hCD;
                    16'hE8E6: data_out = 8'hCE;
                    16'hE8E7: data_out = 8'hCF;
                    16'hE8E8: data_out = 8'hD0;
                    16'hE8E9: data_out = 8'hD1;
                    16'hE8EA: data_out = 8'hD2;
                    16'hE8EB: data_out = 8'hD3;
                    16'hE8EC: data_out = 8'hD4;
                    16'hE8ED: data_out = 8'hD5;
                    16'hE8EE: data_out = 8'hD6;
                    16'hE8EF: data_out = 8'hD7;
                    16'hE8F0: data_out = 8'hD8;
                    16'hE8F1: data_out = 8'hD9;
                    16'hE8F2: data_out = 8'hDA;
                    16'hE8F3: data_out = 8'hDB;
                    16'hE8F4: data_out = 8'hDC;
                    16'hE8F5: data_out = 8'hDD;
                    16'hE8F6: data_out = 8'hDE;
                    16'hE8F7: data_out = 8'hDF;
                    16'hE8F8: data_out = 8'hE0;
                    16'hE8F9: data_out = 8'hE1;
                    16'hE8FA: data_out = 8'hE2;
                    16'hE8FB: data_out = 8'hE3;
                    16'hE8FC: data_out = 8'hE4;
                    16'hE8FD: data_out = 8'hE5;
                    16'hE8FE: data_out = 8'hE6;
                    16'hE8FF: data_out = 8'hE7;
                    16'hE900: data_out = 8'hE9;
                    16'hE901: data_out = 8'hE8;
                    16'hE902: data_out = 8'hE7;
                    16'hE903: data_out = 8'hE6;
                    16'hE904: data_out = 8'hE5;
                    16'hE905: data_out = 8'hE4;
                    16'hE906: data_out = 8'hE3;
                    16'hE907: data_out = 8'hE2;
                    16'hE908: data_out = 8'hE1;
                    16'hE909: data_out = 8'hE0;
                    16'hE90A: data_out = 8'hDF;
                    16'hE90B: data_out = 8'hDE;
                    16'hE90C: data_out = 8'hDD;
                    16'hE90D: data_out = 8'hDC;
                    16'hE90E: data_out = 8'hDB;
                    16'hE90F: data_out = 8'hDA;
                    16'hE910: data_out = 8'hD9;
                    16'hE911: data_out = 8'hD8;
                    16'hE912: data_out = 8'hD7;
                    16'hE913: data_out = 8'hD6;
                    16'hE914: data_out = 8'hD5;
                    16'hE915: data_out = 8'hD4;
                    16'hE916: data_out = 8'hD3;
                    16'hE917: data_out = 8'hD2;
                    16'hE918: data_out = 8'hD1;
                    16'hE919: data_out = 8'hD0;
                    16'hE91A: data_out = 8'hCF;
                    16'hE91B: data_out = 8'hCE;
                    16'hE91C: data_out = 8'hCD;
                    16'hE91D: data_out = 8'hCC;
                    16'hE91E: data_out = 8'hCB;
                    16'hE91F: data_out = 8'hCA;
                    16'hE920: data_out = 8'hC9;
                    16'hE921: data_out = 8'hC8;
                    16'hE922: data_out = 8'hC7;
                    16'hE923: data_out = 8'hC6;
                    16'hE924: data_out = 8'hC5;
                    16'hE925: data_out = 8'hC4;
                    16'hE926: data_out = 8'hC3;
                    16'hE927: data_out = 8'hC2;
                    16'hE928: data_out = 8'hC1;
                    16'hE929: data_out = 8'hC0;
                    16'hE92A: data_out = 8'hBF;
                    16'hE92B: data_out = 8'hBE;
                    16'hE92C: data_out = 8'hBD;
                    16'hE92D: data_out = 8'hBC;
                    16'hE92E: data_out = 8'hBB;
                    16'hE92F: data_out = 8'hBA;
                    16'hE930: data_out = 8'hB9;
                    16'hE931: data_out = 8'hB8;
                    16'hE932: data_out = 8'hB7;
                    16'hE933: data_out = 8'hB6;
                    16'hE934: data_out = 8'hB5;
                    16'hE935: data_out = 8'hB4;
                    16'hE936: data_out = 8'hB3;
                    16'hE937: data_out = 8'hB2;
                    16'hE938: data_out = 8'hB1;
                    16'hE939: data_out = 8'hB0;
                    16'hE93A: data_out = 8'hAF;
                    16'hE93B: data_out = 8'hAE;
                    16'hE93C: data_out = 8'hAD;
                    16'hE93D: data_out = 8'hAC;
                    16'hE93E: data_out = 8'hAB;
                    16'hE93F: data_out = 8'hAA;
                    16'hE940: data_out = 8'hA9;
                    16'hE941: data_out = 8'hA8;
                    16'hE942: data_out = 8'hA7;
                    16'hE943: data_out = 8'hA6;
                    16'hE944: data_out = 8'hA5;
                    16'hE945: data_out = 8'hA4;
                    16'hE946: data_out = 8'hA3;
                    16'hE947: data_out = 8'hA2;
                    16'hE948: data_out = 8'hA1;
                    16'hE949: data_out = 8'hA0;
                    16'hE94A: data_out = 8'h9F;
                    16'hE94B: data_out = 8'h9E;
                    16'hE94C: data_out = 8'h9D;
                    16'hE94D: data_out = 8'h9C;
                    16'hE94E: data_out = 8'h9B;
                    16'hE94F: data_out = 8'h9A;
                    16'hE950: data_out = 8'h99;
                    16'hE951: data_out = 8'h98;
                    16'hE952: data_out = 8'h97;
                    16'hE953: data_out = 8'h96;
                    16'hE954: data_out = 8'h95;
                    16'hE955: data_out = 8'h94;
                    16'hE956: data_out = 8'h93;
                    16'hE957: data_out = 8'h92;
                    16'hE958: data_out = 8'h91;
                    16'hE959: data_out = 8'h90;
                    16'hE95A: data_out = 8'h8F;
                    16'hE95B: data_out = 8'h8E;
                    16'hE95C: data_out = 8'h8D;
                    16'hE95D: data_out = 8'h8C;
                    16'hE95E: data_out = 8'h8B;
                    16'hE95F: data_out = 8'h8A;
                    16'hE960: data_out = 8'h89;
                    16'hE961: data_out = 8'h88;
                    16'hE962: data_out = 8'h87;
                    16'hE963: data_out = 8'h86;
                    16'hE964: data_out = 8'h85;
                    16'hE965: data_out = 8'h84;
                    16'hE966: data_out = 8'h83;
                    16'hE967: data_out = 8'h82;
                    16'hE968: data_out = 8'h81;
                    16'hE969: data_out = 8'h0;
                    16'hE96A: data_out = 8'h1;
                    16'hE96B: data_out = 8'h2;
                    16'hE96C: data_out = 8'h3;
                    16'hE96D: data_out = 8'h4;
                    16'hE96E: data_out = 8'h5;
                    16'hE96F: data_out = 8'h6;
                    16'hE970: data_out = 8'h7;
                    16'hE971: data_out = 8'h8;
                    16'hE972: data_out = 8'h9;
                    16'hE973: data_out = 8'hA;
                    16'hE974: data_out = 8'hB;
                    16'hE975: data_out = 8'hC;
                    16'hE976: data_out = 8'hD;
                    16'hE977: data_out = 8'hE;
                    16'hE978: data_out = 8'hF;
                    16'hE979: data_out = 8'h10;
                    16'hE97A: data_out = 8'h11;
                    16'hE97B: data_out = 8'h12;
                    16'hE97C: data_out = 8'h13;
                    16'hE97D: data_out = 8'h14;
                    16'hE97E: data_out = 8'h15;
                    16'hE97F: data_out = 8'h16;
                    16'hE980: data_out = 8'hE9;
                    16'hE981: data_out = 8'hEA;
                    16'hE982: data_out = 8'hEB;
                    16'hE983: data_out = 8'hEC;
                    16'hE984: data_out = 8'hED;
                    16'hE985: data_out = 8'hEE;
                    16'hE986: data_out = 8'hEF;
                    16'hE987: data_out = 8'hF0;
                    16'hE988: data_out = 8'hF1;
                    16'hE989: data_out = 8'hF2;
                    16'hE98A: data_out = 8'hF3;
                    16'hE98B: data_out = 8'hF4;
                    16'hE98C: data_out = 8'hF5;
                    16'hE98D: data_out = 8'hF6;
                    16'hE98E: data_out = 8'hF7;
                    16'hE98F: data_out = 8'hF8;
                    16'hE990: data_out = 8'hF9;
                    16'hE991: data_out = 8'hFA;
                    16'hE992: data_out = 8'hFB;
                    16'hE993: data_out = 8'hFC;
                    16'hE994: data_out = 8'hFD;
                    16'hE995: data_out = 8'hFE;
                    16'hE996: data_out = 8'hFF;
                    16'hE997: data_out = 8'h80;
                    16'hE998: data_out = 8'h81;
                    16'hE999: data_out = 8'h82;
                    16'hE99A: data_out = 8'h83;
                    16'hE99B: data_out = 8'h84;
                    16'hE99C: data_out = 8'h85;
                    16'hE99D: data_out = 8'h86;
                    16'hE99E: data_out = 8'h87;
                    16'hE99F: data_out = 8'h88;
                    16'hE9A0: data_out = 8'h89;
                    16'hE9A1: data_out = 8'h8A;
                    16'hE9A2: data_out = 8'h8B;
                    16'hE9A3: data_out = 8'h8C;
                    16'hE9A4: data_out = 8'h8D;
                    16'hE9A5: data_out = 8'h8E;
                    16'hE9A6: data_out = 8'h8F;
                    16'hE9A7: data_out = 8'h90;
                    16'hE9A8: data_out = 8'h91;
                    16'hE9A9: data_out = 8'h92;
                    16'hE9AA: data_out = 8'h93;
                    16'hE9AB: data_out = 8'h94;
                    16'hE9AC: data_out = 8'h95;
                    16'hE9AD: data_out = 8'h96;
                    16'hE9AE: data_out = 8'h97;
                    16'hE9AF: data_out = 8'h98;
                    16'hE9B0: data_out = 8'h99;
                    16'hE9B1: data_out = 8'h9A;
                    16'hE9B2: data_out = 8'h9B;
                    16'hE9B3: data_out = 8'h9C;
                    16'hE9B4: data_out = 8'h9D;
                    16'hE9B5: data_out = 8'h9E;
                    16'hE9B6: data_out = 8'h9F;
                    16'hE9B7: data_out = 8'hA0;
                    16'hE9B8: data_out = 8'hA1;
                    16'hE9B9: data_out = 8'hA2;
                    16'hE9BA: data_out = 8'hA3;
                    16'hE9BB: data_out = 8'hA4;
                    16'hE9BC: data_out = 8'hA5;
                    16'hE9BD: data_out = 8'hA6;
                    16'hE9BE: data_out = 8'hA7;
                    16'hE9BF: data_out = 8'hA8;
                    16'hE9C0: data_out = 8'hA9;
                    16'hE9C1: data_out = 8'hAA;
                    16'hE9C2: data_out = 8'hAB;
                    16'hE9C3: data_out = 8'hAC;
                    16'hE9C4: data_out = 8'hAD;
                    16'hE9C5: data_out = 8'hAE;
                    16'hE9C6: data_out = 8'hAF;
                    16'hE9C7: data_out = 8'hB0;
                    16'hE9C8: data_out = 8'hB1;
                    16'hE9C9: data_out = 8'hB2;
                    16'hE9CA: data_out = 8'hB3;
                    16'hE9CB: data_out = 8'hB4;
                    16'hE9CC: data_out = 8'hB5;
                    16'hE9CD: data_out = 8'hB6;
                    16'hE9CE: data_out = 8'hB7;
                    16'hE9CF: data_out = 8'hB8;
                    16'hE9D0: data_out = 8'hB9;
                    16'hE9D1: data_out = 8'hBA;
                    16'hE9D2: data_out = 8'hBB;
                    16'hE9D3: data_out = 8'hBC;
                    16'hE9D4: data_out = 8'hBD;
                    16'hE9D5: data_out = 8'hBE;
                    16'hE9D6: data_out = 8'hBF;
                    16'hE9D7: data_out = 8'hC0;
                    16'hE9D8: data_out = 8'hC1;
                    16'hE9D9: data_out = 8'hC2;
                    16'hE9DA: data_out = 8'hC3;
                    16'hE9DB: data_out = 8'hC4;
                    16'hE9DC: data_out = 8'hC5;
                    16'hE9DD: data_out = 8'hC6;
                    16'hE9DE: data_out = 8'hC7;
                    16'hE9DF: data_out = 8'hC8;
                    16'hE9E0: data_out = 8'hC9;
                    16'hE9E1: data_out = 8'hCA;
                    16'hE9E2: data_out = 8'hCB;
                    16'hE9E3: data_out = 8'hCC;
                    16'hE9E4: data_out = 8'hCD;
                    16'hE9E5: data_out = 8'hCE;
                    16'hE9E6: data_out = 8'hCF;
                    16'hE9E7: data_out = 8'hD0;
                    16'hE9E8: data_out = 8'hD1;
                    16'hE9E9: data_out = 8'hD2;
                    16'hE9EA: data_out = 8'hD3;
                    16'hE9EB: data_out = 8'hD4;
                    16'hE9EC: data_out = 8'hD5;
                    16'hE9ED: data_out = 8'hD6;
                    16'hE9EE: data_out = 8'hD7;
                    16'hE9EF: data_out = 8'hD8;
                    16'hE9F0: data_out = 8'hD9;
                    16'hE9F1: data_out = 8'hDA;
                    16'hE9F2: data_out = 8'hDB;
                    16'hE9F3: data_out = 8'hDC;
                    16'hE9F4: data_out = 8'hDD;
                    16'hE9F5: data_out = 8'hDE;
                    16'hE9F6: data_out = 8'hDF;
                    16'hE9F7: data_out = 8'hE0;
                    16'hE9F8: data_out = 8'hE1;
                    16'hE9F9: data_out = 8'hE2;
                    16'hE9FA: data_out = 8'hE3;
                    16'hE9FB: data_out = 8'hE4;
                    16'hE9FC: data_out = 8'hE5;
                    16'hE9FD: data_out = 8'hE6;
                    16'hE9FE: data_out = 8'hE7;
                    16'hE9FF: data_out = 8'hE8;
                    16'hEA00: data_out = 8'hEA;
                    16'hEA01: data_out = 8'hE9;
                    16'hEA02: data_out = 8'hE8;
                    16'hEA03: data_out = 8'hE7;
                    16'hEA04: data_out = 8'hE6;
                    16'hEA05: data_out = 8'hE5;
                    16'hEA06: data_out = 8'hE4;
                    16'hEA07: data_out = 8'hE3;
                    16'hEA08: data_out = 8'hE2;
                    16'hEA09: data_out = 8'hE1;
                    16'hEA0A: data_out = 8'hE0;
                    16'hEA0B: data_out = 8'hDF;
                    16'hEA0C: data_out = 8'hDE;
                    16'hEA0D: data_out = 8'hDD;
                    16'hEA0E: data_out = 8'hDC;
                    16'hEA0F: data_out = 8'hDB;
                    16'hEA10: data_out = 8'hDA;
                    16'hEA11: data_out = 8'hD9;
                    16'hEA12: data_out = 8'hD8;
                    16'hEA13: data_out = 8'hD7;
                    16'hEA14: data_out = 8'hD6;
                    16'hEA15: data_out = 8'hD5;
                    16'hEA16: data_out = 8'hD4;
                    16'hEA17: data_out = 8'hD3;
                    16'hEA18: data_out = 8'hD2;
                    16'hEA19: data_out = 8'hD1;
                    16'hEA1A: data_out = 8'hD0;
                    16'hEA1B: data_out = 8'hCF;
                    16'hEA1C: data_out = 8'hCE;
                    16'hEA1D: data_out = 8'hCD;
                    16'hEA1E: data_out = 8'hCC;
                    16'hEA1F: data_out = 8'hCB;
                    16'hEA20: data_out = 8'hCA;
                    16'hEA21: data_out = 8'hC9;
                    16'hEA22: data_out = 8'hC8;
                    16'hEA23: data_out = 8'hC7;
                    16'hEA24: data_out = 8'hC6;
                    16'hEA25: data_out = 8'hC5;
                    16'hEA26: data_out = 8'hC4;
                    16'hEA27: data_out = 8'hC3;
                    16'hEA28: data_out = 8'hC2;
                    16'hEA29: data_out = 8'hC1;
                    16'hEA2A: data_out = 8'hC0;
                    16'hEA2B: data_out = 8'hBF;
                    16'hEA2C: data_out = 8'hBE;
                    16'hEA2D: data_out = 8'hBD;
                    16'hEA2E: data_out = 8'hBC;
                    16'hEA2F: data_out = 8'hBB;
                    16'hEA30: data_out = 8'hBA;
                    16'hEA31: data_out = 8'hB9;
                    16'hEA32: data_out = 8'hB8;
                    16'hEA33: data_out = 8'hB7;
                    16'hEA34: data_out = 8'hB6;
                    16'hEA35: data_out = 8'hB5;
                    16'hEA36: data_out = 8'hB4;
                    16'hEA37: data_out = 8'hB3;
                    16'hEA38: data_out = 8'hB2;
                    16'hEA39: data_out = 8'hB1;
                    16'hEA3A: data_out = 8'hB0;
                    16'hEA3B: data_out = 8'hAF;
                    16'hEA3C: data_out = 8'hAE;
                    16'hEA3D: data_out = 8'hAD;
                    16'hEA3E: data_out = 8'hAC;
                    16'hEA3F: data_out = 8'hAB;
                    16'hEA40: data_out = 8'hAA;
                    16'hEA41: data_out = 8'hA9;
                    16'hEA42: data_out = 8'hA8;
                    16'hEA43: data_out = 8'hA7;
                    16'hEA44: data_out = 8'hA6;
                    16'hEA45: data_out = 8'hA5;
                    16'hEA46: data_out = 8'hA4;
                    16'hEA47: data_out = 8'hA3;
                    16'hEA48: data_out = 8'hA2;
                    16'hEA49: data_out = 8'hA1;
                    16'hEA4A: data_out = 8'hA0;
                    16'hEA4B: data_out = 8'h9F;
                    16'hEA4C: data_out = 8'h9E;
                    16'hEA4D: data_out = 8'h9D;
                    16'hEA4E: data_out = 8'h9C;
                    16'hEA4F: data_out = 8'h9B;
                    16'hEA50: data_out = 8'h9A;
                    16'hEA51: data_out = 8'h99;
                    16'hEA52: data_out = 8'h98;
                    16'hEA53: data_out = 8'h97;
                    16'hEA54: data_out = 8'h96;
                    16'hEA55: data_out = 8'h95;
                    16'hEA56: data_out = 8'h94;
                    16'hEA57: data_out = 8'h93;
                    16'hEA58: data_out = 8'h92;
                    16'hEA59: data_out = 8'h91;
                    16'hEA5A: data_out = 8'h90;
                    16'hEA5B: data_out = 8'h8F;
                    16'hEA5C: data_out = 8'h8E;
                    16'hEA5D: data_out = 8'h8D;
                    16'hEA5E: data_out = 8'h8C;
                    16'hEA5F: data_out = 8'h8B;
                    16'hEA60: data_out = 8'h8A;
                    16'hEA61: data_out = 8'h89;
                    16'hEA62: data_out = 8'h88;
                    16'hEA63: data_out = 8'h87;
                    16'hEA64: data_out = 8'h86;
                    16'hEA65: data_out = 8'h85;
                    16'hEA66: data_out = 8'h84;
                    16'hEA67: data_out = 8'h83;
                    16'hEA68: data_out = 8'h82;
                    16'hEA69: data_out = 8'h81;
                    16'hEA6A: data_out = 8'h0;
                    16'hEA6B: data_out = 8'h1;
                    16'hEA6C: data_out = 8'h2;
                    16'hEA6D: data_out = 8'h3;
                    16'hEA6E: data_out = 8'h4;
                    16'hEA6F: data_out = 8'h5;
                    16'hEA70: data_out = 8'h6;
                    16'hEA71: data_out = 8'h7;
                    16'hEA72: data_out = 8'h8;
                    16'hEA73: data_out = 8'h9;
                    16'hEA74: data_out = 8'hA;
                    16'hEA75: data_out = 8'hB;
                    16'hEA76: data_out = 8'hC;
                    16'hEA77: data_out = 8'hD;
                    16'hEA78: data_out = 8'hE;
                    16'hEA79: data_out = 8'hF;
                    16'hEA7A: data_out = 8'h10;
                    16'hEA7B: data_out = 8'h11;
                    16'hEA7C: data_out = 8'h12;
                    16'hEA7D: data_out = 8'h13;
                    16'hEA7E: data_out = 8'h14;
                    16'hEA7F: data_out = 8'h15;
                    16'hEA80: data_out = 8'hEA;
                    16'hEA81: data_out = 8'hEB;
                    16'hEA82: data_out = 8'hEC;
                    16'hEA83: data_out = 8'hED;
                    16'hEA84: data_out = 8'hEE;
                    16'hEA85: data_out = 8'hEF;
                    16'hEA86: data_out = 8'hF0;
                    16'hEA87: data_out = 8'hF1;
                    16'hEA88: data_out = 8'hF2;
                    16'hEA89: data_out = 8'hF3;
                    16'hEA8A: data_out = 8'hF4;
                    16'hEA8B: data_out = 8'hF5;
                    16'hEA8C: data_out = 8'hF6;
                    16'hEA8D: data_out = 8'hF7;
                    16'hEA8E: data_out = 8'hF8;
                    16'hEA8F: data_out = 8'hF9;
                    16'hEA90: data_out = 8'hFA;
                    16'hEA91: data_out = 8'hFB;
                    16'hEA92: data_out = 8'hFC;
                    16'hEA93: data_out = 8'hFD;
                    16'hEA94: data_out = 8'hFE;
                    16'hEA95: data_out = 8'hFF;
                    16'hEA96: data_out = 8'h80;
                    16'hEA97: data_out = 8'h81;
                    16'hEA98: data_out = 8'h82;
                    16'hEA99: data_out = 8'h83;
                    16'hEA9A: data_out = 8'h84;
                    16'hEA9B: data_out = 8'h85;
                    16'hEA9C: data_out = 8'h86;
                    16'hEA9D: data_out = 8'h87;
                    16'hEA9E: data_out = 8'h88;
                    16'hEA9F: data_out = 8'h89;
                    16'hEAA0: data_out = 8'h8A;
                    16'hEAA1: data_out = 8'h8B;
                    16'hEAA2: data_out = 8'h8C;
                    16'hEAA3: data_out = 8'h8D;
                    16'hEAA4: data_out = 8'h8E;
                    16'hEAA5: data_out = 8'h8F;
                    16'hEAA6: data_out = 8'h90;
                    16'hEAA7: data_out = 8'h91;
                    16'hEAA8: data_out = 8'h92;
                    16'hEAA9: data_out = 8'h93;
                    16'hEAAA: data_out = 8'h94;
                    16'hEAAB: data_out = 8'h95;
                    16'hEAAC: data_out = 8'h96;
                    16'hEAAD: data_out = 8'h97;
                    16'hEAAE: data_out = 8'h98;
                    16'hEAAF: data_out = 8'h99;
                    16'hEAB0: data_out = 8'h9A;
                    16'hEAB1: data_out = 8'h9B;
                    16'hEAB2: data_out = 8'h9C;
                    16'hEAB3: data_out = 8'h9D;
                    16'hEAB4: data_out = 8'h9E;
                    16'hEAB5: data_out = 8'h9F;
                    16'hEAB6: data_out = 8'hA0;
                    16'hEAB7: data_out = 8'hA1;
                    16'hEAB8: data_out = 8'hA2;
                    16'hEAB9: data_out = 8'hA3;
                    16'hEABA: data_out = 8'hA4;
                    16'hEABB: data_out = 8'hA5;
                    16'hEABC: data_out = 8'hA6;
                    16'hEABD: data_out = 8'hA7;
                    16'hEABE: data_out = 8'hA8;
                    16'hEABF: data_out = 8'hA9;
                    16'hEAC0: data_out = 8'hAA;
                    16'hEAC1: data_out = 8'hAB;
                    16'hEAC2: data_out = 8'hAC;
                    16'hEAC3: data_out = 8'hAD;
                    16'hEAC4: data_out = 8'hAE;
                    16'hEAC5: data_out = 8'hAF;
                    16'hEAC6: data_out = 8'hB0;
                    16'hEAC7: data_out = 8'hB1;
                    16'hEAC8: data_out = 8'hB2;
                    16'hEAC9: data_out = 8'hB3;
                    16'hEACA: data_out = 8'hB4;
                    16'hEACB: data_out = 8'hB5;
                    16'hEACC: data_out = 8'hB6;
                    16'hEACD: data_out = 8'hB7;
                    16'hEACE: data_out = 8'hB8;
                    16'hEACF: data_out = 8'hB9;
                    16'hEAD0: data_out = 8'hBA;
                    16'hEAD1: data_out = 8'hBB;
                    16'hEAD2: data_out = 8'hBC;
                    16'hEAD3: data_out = 8'hBD;
                    16'hEAD4: data_out = 8'hBE;
                    16'hEAD5: data_out = 8'hBF;
                    16'hEAD6: data_out = 8'hC0;
                    16'hEAD7: data_out = 8'hC1;
                    16'hEAD8: data_out = 8'hC2;
                    16'hEAD9: data_out = 8'hC3;
                    16'hEADA: data_out = 8'hC4;
                    16'hEADB: data_out = 8'hC5;
                    16'hEADC: data_out = 8'hC6;
                    16'hEADD: data_out = 8'hC7;
                    16'hEADE: data_out = 8'hC8;
                    16'hEADF: data_out = 8'hC9;
                    16'hEAE0: data_out = 8'hCA;
                    16'hEAE1: data_out = 8'hCB;
                    16'hEAE2: data_out = 8'hCC;
                    16'hEAE3: data_out = 8'hCD;
                    16'hEAE4: data_out = 8'hCE;
                    16'hEAE5: data_out = 8'hCF;
                    16'hEAE6: data_out = 8'hD0;
                    16'hEAE7: data_out = 8'hD1;
                    16'hEAE8: data_out = 8'hD2;
                    16'hEAE9: data_out = 8'hD3;
                    16'hEAEA: data_out = 8'hD4;
                    16'hEAEB: data_out = 8'hD5;
                    16'hEAEC: data_out = 8'hD6;
                    16'hEAED: data_out = 8'hD7;
                    16'hEAEE: data_out = 8'hD8;
                    16'hEAEF: data_out = 8'hD9;
                    16'hEAF0: data_out = 8'hDA;
                    16'hEAF1: data_out = 8'hDB;
                    16'hEAF2: data_out = 8'hDC;
                    16'hEAF3: data_out = 8'hDD;
                    16'hEAF4: data_out = 8'hDE;
                    16'hEAF5: data_out = 8'hDF;
                    16'hEAF6: data_out = 8'hE0;
                    16'hEAF7: data_out = 8'hE1;
                    16'hEAF8: data_out = 8'hE2;
                    16'hEAF9: data_out = 8'hE3;
                    16'hEAFA: data_out = 8'hE4;
                    16'hEAFB: data_out = 8'hE5;
                    16'hEAFC: data_out = 8'hE6;
                    16'hEAFD: data_out = 8'hE7;
                    16'hEAFE: data_out = 8'hE8;
                    16'hEAFF: data_out = 8'hE9;
                    16'hEB00: data_out = 8'hEB;
                    16'hEB01: data_out = 8'hEA;
                    16'hEB02: data_out = 8'hE9;
                    16'hEB03: data_out = 8'hE8;
                    16'hEB04: data_out = 8'hE7;
                    16'hEB05: data_out = 8'hE6;
                    16'hEB06: data_out = 8'hE5;
                    16'hEB07: data_out = 8'hE4;
                    16'hEB08: data_out = 8'hE3;
                    16'hEB09: data_out = 8'hE2;
                    16'hEB0A: data_out = 8'hE1;
                    16'hEB0B: data_out = 8'hE0;
                    16'hEB0C: data_out = 8'hDF;
                    16'hEB0D: data_out = 8'hDE;
                    16'hEB0E: data_out = 8'hDD;
                    16'hEB0F: data_out = 8'hDC;
                    16'hEB10: data_out = 8'hDB;
                    16'hEB11: data_out = 8'hDA;
                    16'hEB12: data_out = 8'hD9;
                    16'hEB13: data_out = 8'hD8;
                    16'hEB14: data_out = 8'hD7;
                    16'hEB15: data_out = 8'hD6;
                    16'hEB16: data_out = 8'hD5;
                    16'hEB17: data_out = 8'hD4;
                    16'hEB18: data_out = 8'hD3;
                    16'hEB19: data_out = 8'hD2;
                    16'hEB1A: data_out = 8'hD1;
                    16'hEB1B: data_out = 8'hD0;
                    16'hEB1C: data_out = 8'hCF;
                    16'hEB1D: data_out = 8'hCE;
                    16'hEB1E: data_out = 8'hCD;
                    16'hEB1F: data_out = 8'hCC;
                    16'hEB20: data_out = 8'hCB;
                    16'hEB21: data_out = 8'hCA;
                    16'hEB22: data_out = 8'hC9;
                    16'hEB23: data_out = 8'hC8;
                    16'hEB24: data_out = 8'hC7;
                    16'hEB25: data_out = 8'hC6;
                    16'hEB26: data_out = 8'hC5;
                    16'hEB27: data_out = 8'hC4;
                    16'hEB28: data_out = 8'hC3;
                    16'hEB29: data_out = 8'hC2;
                    16'hEB2A: data_out = 8'hC1;
                    16'hEB2B: data_out = 8'hC0;
                    16'hEB2C: data_out = 8'hBF;
                    16'hEB2D: data_out = 8'hBE;
                    16'hEB2E: data_out = 8'hBD;
                    16'hEB2F: data_out = 8'hBC;
                    16'hEB30: data_out = 8'hBB;
                    16'hEB31: data_out = 8'hBA;
                    16'hEB32: data_out = 8'hB9;
                    16'hEB33: data_out = 8'hB8;
                    16'hEB34: data_out = 8'hB7;
                    16'hEB35: data_out = 8'hB6;
                    16'hEB36: data_out = 8'hB5;
                    16'hEB37: data_out = 8'hB4;
                    16'hEB38: data_out = 8'hB3;
                    16'hEB39: data_out = 8'hB2;
                    16'hEB3A: data_out = 8'hB1;
                    16'hEB3B: data_out = 8'hB0;
                    16'hEB3C: data_out = 8'hAF;
                    16'hEB3D: data_out = 8'hAE;
                    16'hEB3E: data_out = 8'hAD;
                    16'hEB3F: data_out = 8'hAC;
                    16'hEB40: data_out = 8'hAB;
                    16'hEB41: data_out = 8'hAA;
                    16'hEB42: data_out = 8'hA9;
                    16'hEB43: data_out = 8'hA8;
                    16'hEB44: data_out = 8'hA7;
                    16'hEB45: data_out = 8'hA6;
                    16'hEB46: data_out = 8'hA5;
                    16'hEB47: data_out = 8'hA4;
                    16'hEB48: data_out = 8'hA3;
                    16'hEB49: data_out = 8'hA2;
                    16'hEB4A: data_out = 8'hA1;
                    16'hEB4B: data_out = 8'hA0;
                    16'hEB4C: data_out = 8'h9F;
                    16'hEB4D: data_out = 8'h9E;
                    16'hEB4E: data_out = 8'h9D;
                    16'hEB4F: data_out = 8'h9C;
                    16'hEB50: data_out = 8'h9B;
                    16'hEB51: data_out = 8'h9A;
                    16'hEB52: data_out = 8'h99;
                    16'hEB53: data_out = 8'h98;
                    16'hEB54: data_out = 8'h97;
                    16'hEB55: data_out = 8'h96;
                    16'hEB56: data_out = 8'h95;
                    16'hEB57: data_out = 8'h94;
                    16'hEB58: data_out = 8'h93;
                    16'hEB59: data_out = 8'h92;
                    16'hEB5A: data_out = 8'h91;
                    16'hEB5B: data_out = 8'h90;
                    16'hEB5C: data_out = 8'h8F;
                    16'hEB5D: data_out = 8'h8E;
                    16'hEB5E: data_out = 8'h8D;
                    16'hEB5F: data_out = 8'h8C;
                    16'hEB60: data_out = 8'h8B;
                    16'hEB61: data_out = 8'h8A;
                    16'hEB62: data_out = 8'h89;
                    16'hEB63: data_out = 8'h88;
                    16'hEB64: data_out = 8'h87;
                    16'hEB65: data_out = 8'h86;
                    16'hEB66: data_out = 8'h85;
                    16'hEB67: data_out = 8'h84;
                    16'hEB68: data_out = 8'h83;
                    16'hEB69: data_out = 8'h82;
                    16'hEB6A: data_out = 8'h81;
                    16'hEB6B: data_out = 8'h0;
                    16'hEB6C: data_out = 8'h1;
                    16'hEB6D: data_out = 8'h2;
                    16'hEB6E: data_out = 8'h3;
                    16'hEB6F: data_out = 8'h4;
                    16'hEB70: data_out = 8'h5;
                    16'hEB71: data_out = 8'h6;
                    16'hEB72: data_out = 8'h7;
                    16'hEB73: data_out = 8'h8;
                    16'hEB74: data_out = 8'h9;
                    16'hEB75: data_out = 8'hA;
                    16'hEB76: data_out = 8'hB;
                    16'hEB77: data_out = 8'hC;
                    16'hEB78: data_out = 8'hD;
                    16'hEB79: data_out = 8'hE;
                    16'hEB7A: data_out = 8'hF;
                    16'hEB7B: data_out = 8'h10;
                    16'hEB7C: data_out = 8'h11;
                    16'hEB7D: data_out = 8'h12;
                    16'hEB7E: data_out = 8'h13;
                    16'hEB7F: data_out = 8'h14;
                    16'hEB80: data_out = 8'hEB;
                    16'hEB81: data_out = 8'hEC;
                    16'hEB82: data_out = 8'hED;
                    16'hEB83: data_out = 8'hEE;
                    16'hEB84: data_out = 8'hEF;
                    16'hEB85: data_out = 8'hF0;
                    16'hEB86: data_out = 8'hF1;
                    16'hEB87: data_out = 8'hF2;
                    16'hEB88: data_out = 8'hF3;
                    16'hEB89: data_out = 8'hF4;
                    16'hEB8A: data_out = 8'hF5;
                    16'hEB8B: data_out = 8'hF6;
                    16'hEB8C: data_out = 8'hF7;
                    16'hEB8D: data_out = 8'hF8;
                    16'hEB8E: data_out = 8'hF9;
                    16'hEB8F: data_out = 8'hFA;
                    16'hEB90: data_out = 8'hFB;
                    16'hEB91: data_out = 8'hFC;
                    16'hEB92: data_out = 8'hFD;
                    16'hEB93: data_out = 8'hFE;
                    16'hEB94: data_out = 8'hFF;
                    16'hEB95: data_out = 8'h80;
                    16'hEB96: data_out = 8'h81;
                    16'hEB97: data_out = 8'h82;
                    16'hEB98: data_out = 8'h83;
                    16'hEB99: data_out = 8'h84;
                    16'hEB9A: data_out = 8'h85;
                    16'hEB9B: data_out = 8'h86;
                    16'hEB9C: data_out = 8'h87;
                    16'hEB9D: data_out = 8'h88;
                    16'hEB9E: data_out = 8'h89;
                    16'hEB9F: data_out = 8'h8A;
                    16'hEBA0: data_out = 8'h8B;
                    16'hEBA1: data_out = 8'h8C;
                    16'hEBA2: data_out = 8'h8D;
                    16'hEBA3: data_out = 8'h8E;
                    16'hEBA4: data_out = 8'h8F;
                    16'hEBA5: data_out = 8'h90;
                    16'hEBA6: data_out = 8'h91;
                    16'hEBA7: data_out = 8'h92;
                    16'hEBA8: data_out = 8'h93;
                    16'hEBA9: data_out = 8'h94;
                    16'hEBAA: data_out = 8'h95;
                    16'hEBAB: data_out = 8'h96;
                    16'hEBAC: data_out = 8'h97;
                    16'hEBAD: data_out = 8'h98;
                    16'hEBAE: data_out = 8'h99;
                    16'hEBAF: data_out = 8'h9A;
                    16'hEBB0: data_out = 8'h9B;
                    16'hEBB1: data_out = 8'h9C;
                    16'hEBB2: data_out = 8'h9D;
                    16'hEBB3: data_out = 8'h9E;
                    16'hEBB4: data_out = 8'h9F;
                    16'hEBB5: data_out = 8'hA0;
                    16'hEBB6: data_out = 8'hA1;
                    16'hEBB7: data_out = 8'hA2;
                    16'hEBB8: data_out = 8'hA3;
                    16'hEBB9: data_out = 8'hA4;
                    16'hEBBA: data_out = 8'hA5;
                    16'hEBBB: data_out = 8'hA6;
                    16'hEBBC: data_out = 8'hA7;
                    16'hEBBD: data_out = 8'hA8;
                    16'hEBBE: data_out = 8'hA9;
                    16'hEBBF: data_out = 8'hAA;
                    16'hEBC0: data_out = 8'hAB;
                    16'hEBC1: data_out = 8'hAC;
                    16'hEBC2: data_out = 8'hAD;
                    16'hEBC3: data_out = 8'hAE;
                    16'hEBC4: data_out = 8'hAF;
                    16'hEBC5: data_out = 8'hB0;
                    16'hEBC6: data_out = 8'hB1;
                    16'hEBC7: data_out = 8'hB2;
                    16'hEBC8: data_out = 8'hB3;
                    16'hEBC9: data_out = 8'hB4;
                    16'hEBCA: data_out = 8'hB5;
                    16'hEBCB: data_out = 8'hB6;
                    16'hEBCC: data_out = 8'hB7;
                    16'hEBCD: data_out = 8'hB8;
                    16'hEBCE: data_out = 8'hB9;
                    16'hEBCF: data_out = 8'hBA;
                    16'hEBD0: data_out = 8'hBB;
                    16'hEBD1: data_out = 8'hBC;
                    16'hEBD2: data_out = 8'hBD;
                    16'hEBD3: data_out = 8'hBE;
                    16'hEBD4: data_out = 8'hBF;
                    16'hEBD5: data_out = 8'hC0;
                    16'hEBD6: data_out = 8'hC1;
                    16'hEBD7: data_out = 8'hC2;
                    16'hEBD8: data_out = 8'hC3;
                    16'hEBD9: data_out = 8'hC4;
                    16'hEBDA: data_out = 8'hC5;
                    16'hEBDB: data_out = 8'hC6;
                    16'hEBDC: data_out = 8'hC7;
                    16'hEBDD: data_out = 8'hC8;
                    16'hEBDE: data_out = 8'hC9;
                    16'hEBDF: data_out = 8'hCA;
                    16'hEBE0: data_out = 8'hCB;
                    16'hEBE1: data_out = 8'hCC;
                    16'hEBE2: data_out = 8'hCD;
                    16'hEBE3: data_out = 8'hCE;
                    16'hEBE4: data_out = 8'hCF;
                    16'hEBE5: data_out = 8'hD0;
                    16'hEBE6: data_out = 8'hD1;
                    16'hEBE7: data_out = 8'hD2;
                    16'hEBE8: data_out = 8'hD3;
                    16'hEBE9: data_out = 8'hD4;
                    16'hEBEA: data_out = 8'hD5;
                    16'hEBEB: data_out = 8'hD6;
                    16'hEBEC: data_out = 8'hD7;
                    16'hEBED: data_out = 8'hD8;
                    16'hEBEE: data_out = 8'hD9;
                    16'hEBEF: data_out = 8'hDA;
                    16'hEBF0: data_out = 8'hDB;
                    16'hEBF1: data_out = 8'hDC;
                    16'hEBF2: data_out = 8'hDD;
                    16'hEBF3: data_out = 8'hDE;
                    16'hEBF4: data_out = 8'hDF;
                    16'hEBF5: data_out = 8'hE0;
                    16'hEBF6: data_out = 8'hE1;
                    16'hEBF7: data_out = 8'hE2;
                    16'hEBF8: data_out = 8'hE3;
                    16'hEBF9: data_out = 8'hE4;
                    16'hEBFA: data_out = 8'hE5;
                    16'hEBFB: data_out = 8'hE6;
                    16'hEBFC: data_out = 8'hE7;
                    16'hEBFD: data_out = 8'hE8;
                    16'hEBFE: data_out = 8'hE9;
                    16'hEBFF: data_out = 8'hEA;
                    16'hEC00: data_out = 8'hEC;
                    16'hEC01: data_out = 8'hEB;
                    16'hEC02: data_out = 8'hEA;
                    16'hEC03: data_out = 8'hE9;
                    16'hEC04: data_out = 8'hE8;
                    16'hEC05: data_out = 8'hE7;
                    16'hEC06: data_out = 8'hE6;
                    16'hEC07: data_out = 8'hE5;
                    16'hEC08: data_out = 8'hE4;
                    16'hEC09: data_out = 8'hE3;
                    16'hEC0A: data_out = 8'hE2;
                    16'hEC0B: data_out = 8'hE1;
                    16'hEC0C: data_out = 8'hE0;
                    16'hEC0D: data_out = 8'hDF;
                    16'hEC0E: data_out = 8'hDE;
                    16'hEC0F: data_out = 8'hDD;
                    16'hEC10: data_out = 8'hDC;
                    16'hEC11: data_out = 8'hDB;
                    16'hEC12: data_out = 8'hDA;
                    16'hEC13: data_out = 8'hD9;
                    16'hEC14: data_out = 8'hD8;
                    16'hEC15: data_out = 8'hD7;
                    16'hEC16: data_out = 8'hD6;
                    16'hEC17: data_out = 8'hD5;
                    16'hEC18: data_out = 8'hD4;
                    16'hEC19: data_out = 8'hD3;
                    16'hEC1A: data_out = 8'hD2;
                    16'hEC1B: data_out = 8'hD1;
                    16'hEC1C: data_out = 8'hD0;
                    16'hEC1D: data_out = 8'hCF;
                    16'hEC1E: data_out = 8'hCE;
                    16'hEC1F: data_out = 8'hCD;
                    16'hEC20: data_out = 8'hCC;
                    16'hEC21: data_out = 8'hCB;
                    16'hEC22: data_out = 8'hCA;
                    16'hEC23: data_out = 8'hC9;
                    16'hEC24: data_out = 8'hC8;
                    16'hEC25: data_out = 8'hC7;
                    16'hEC26: data_out = 8'hC6;
                    16'hEC27: data_out = 8'hC5;
                    16'hEC28: data_out = 8'hC4;
                    16'hEC29: data_out = 8'hC3;
                    16'hEC2A: data_out = 8'hC2;
                    16'hEC2B: data_out = 8'hC1;
                    16'hEC2C: data_out = 8'hC0;
                    16'hEC2D: data_out = 8'hBF;
                    16'hEC2E: data_out = 8'hBE;
                    16'hEC2F: data_out = 8'hBD;
                    16'hEC30: data_out = 8'hBC;
                    16'hEC31: data_out = 8'hBB;
                    16'hEC32: data_out = 8'hBA;
                    16'hEC33: data_out = 8'hB9;
                    16'hEC34: data_out = 8'hB8;
                    16'hEC35: data_out = 8'hB7;
                    16'hEC36: data_out = 8'hB6;
                    16'hEC37: data_out = 8'hB5;
                    16'hEC38: data_out = 8'hB4;
                    16'hEC39: data_out = 8'hB3;
                    16'hEC3A: data_out = 8'hB2;
                    16'hEC3B: data_out = 8'hB1;
                    16'hEC3C: data_out = 8'hB0;
                    16'hEC3D: data_out = 8'hAF;
                    16'hEC3E: data_out = 8'hAE;
                    16'hEC3F: data_out = 8'hAD;
                    16'hEC40: data_out = 8'hAC;
                    16'hEC41: data_out = 8'hAB;
                    16'hEC42: data_out = 8'hAA;
                    16'hEC43: data_out = 8'hA9;
                    16'hEC44: data_out = 8'hA8;
                    16'hEC45: data_out = 8'hA7;
                    16'hEC46: data_out = 8'hA6;
                    16'hEC47: data_out = 8'hA5;
                    16'hEC48: data_out = 8'hA4;
                    16'hEC49: data_out = 8'hA3;
                    16'hEC4A: data_out = 8'hA2;
                    16'hEC4B: data_out = 8'hA1;
                    16'hEC4C: data_out = 8'hA0;
                    16'hEC4D: data_out = 8'h9F;
                    16'hEC4E: data_out = 8'h9E;
                    16'hEC4F: data_out = 8'h9D;
                    16'hEC50: data_out = 8'h9C;
                    16'hEC51: data_out = 8'h9B;
                    16'hEC52: data_out = 8'h9A;
                    16'hEC53: data_out = 8'h99;
                    16'hEC54: data_out = 8'h98;
                    16'hEC55: data_out = 8'h97;
                    16'hEC56: data_out = 8'h96;
                    16'hEC57: data_out = 8'h95;
                    16'hEC58: data_out = 8'h94;
                    16'hEC59: data_out = 8'h93;
                    16'hEC5A: data_out = 8'h92;
                    16'hEC5B: data_out = 8'h91;
                    16'hEC5C: data_out = 8'h90;
                    16'hEC5D: data_out = 8'h8F;
                    16'hEC5E: data_out = 8'h8E;
                    16'hEC5F: data_out = 8'h8D;
                    16'hEC60: data_out = 8'h8C;
                    16'hEC61: data_out = 8'h8B;
                    16'hEC62: data_out = 8'h8A;
                    16'hEC63: data_out = 8'h89;
                    16'hEC64: data_out = 8'h88;
                    16'hEC65: data_out = 8'h87;
                    16'hEC66: data_out = 8'h86;
                    16'hEC67: data_out = 8'h85;
                    16'hEC68: data_out = 8'h84;
                    16'hEC69: data_out = 8'h83;
                    16'hEC6A: data_out = 8'h82;
                    16'hEC6B: data_out = 8'h81;
                    16'hEC6C: data_out = 8'h0;
                    16'hEC6D: data_out = 8'h1;
                    16'hEC6E: data_out = 8'h2;
                    16'hEC6F: data_out = 8'h3;
                    16'hEC70: data_out = 8'h4;
                    16'hEC71: data_out = 8'h5;
                    16'hEC72: data_out = 8'h6;
                    16'hEC73: data_out = 8'h7;
                    16'hEC74: data_out = 8'h8;
                    16'hEC75: data_out = 8'h9;
                    16'hEC76: data_out = 8'hA;
                    16'hEC77: data_out = 8'hB;
                    16'hEC78: data_out = 8'hC;
                    16'hEC79: data_out = 8'hD;
                    16'hEC7A: data_out = 8'hE;
                    16'hEC7B: data_out = 8'hF;
                    16'hEC7C: data_out = 8'h10;
                    16'hEC7D: data_out = 8'h11;
                    16'hEC7E: data_out = 8'h12;
                    16'hEC7F: data_out = 8'h13;
                    16'hEC80: data_out = 8'hEC;
                    16'hEC81: data_out = 8'hED;
                    16'hEC82: data_out = 8'hEE;
                    16'hEC83: data_out = 8'hEF;
                    16'hEC84: data_out = 8'hF0;
                    16'hEC85: data_out = 8'hF1;
                    16'hEC86: data_out = 8'hF2;
                    16'hEC87: data_out = 8'hF3;
                    16'hEC88: data_out = 8'hF4;
                    16'hEC89: data_out = 8'hF5;
                    16'hEC8A: data_out = 8'hF6;
                    16'hEC8B: data_out = 8'hF7;
                    16'hEC8C: data_out = 8'hF8;
                    16'hEC8D: data_out = 8'hF9;
                    16'hEC8E: data_out = 8'hFA;
                    16'hEC8F: data_out = 8'hFB;
                    16'hEC90: data_out = 8'hFC;
                    16'hEC91: data_out = 8'hFD;
                    16'hEC92: data_out = 8'hFE;
                    16'hEC93: data_out = 8'hFF;
                    16'hEC94: data_out = 8'h80;
                    16'hEC95: data_out = 8'h81;
                    16'hEC96: data_out = 8'h82;
                    16'hEC97: data_out = 8'h83;
                    16'hEC98: data_out = 8'h84;
                    16'hEC99: data_out = 8'h85;
                    16'hEC9A: data_out = 8'h86;
                    16'hEC9B: data_out = 8'h87;
                    16'hEC9C: data_out = 8'h88;
                    16'hEC9D: data_out = 8'h89;
                    16'hEC9E: data_out = 8'h8A;
                    16'hEC9F: data_out = 8'h8B;
                    16'hECA0: data_out = 8'h8C;
                    16'hECA1: data_out = 8'h8D;
                    16'hECA2: data_out = 8'h8E;
                    16'hECA3: data_out = 8'h8F;
                    16'hECA4: data_out = 8'h90;
                    16'hECA5: data_out = 8'h91;
                    16'hECA6: data_out = 8'h92;
                    16'hECA7: data_out = 8'h93;
                    16'hECA8: data_out = 8'h94;
                    16'hECA9: data_out = 8'h95;
                    16'hECAA: data_out = 8'h96;
                    16'hECAB: data_out = 8'h97;
                    16'hECAC: data_out = 8'h98;
                    16'hECAD: data_out = 8'h99;
                    16'hECAE: data_out = 8'h9A;
                    16'hECAF: data_out = 8'h9B;
                    16'hECB0: data_out = 8'h9C;
                    16'hECB1: data_out = 8'h9D;
                    16'hECB2: data_out = 8'h9E;
                    16'hECB3: data_out = 8'h9F;
                    16'hECB4: data_out = 8'hA0;
                    16'hECB5: data_out = 8'hA1;
                    16'hECB6: data_out = 8'hA2;
                    16'hECB7: data_out = 8'hA3;
                    16'hECB8: data_out = 8'hA4;
                    16'hECB9: data_out = 8'hA5;
                    16'hECBA: data_out = 8'hA6;
                    16'hECBB: data_out = 8'hA7;
                    16'hECBC: data_out = 8'hA8;
                    16'hECBD: data_out = 8'hA9;
                    16'hECBE: data_out = 8'hAA;
                    16'hECBF: data_out = 8'hAB;
                    16'hECC0: data_out = 8'hAC;
                    16'hECC1: data_out = 8'hAD;
                    16'hECC2: data_out = 8'hAE;
                    16'hECC3: data_out = 8'hAF;
                    16'hECC4: data_out = 8'hB0;
                    16'hECC5: data_out = 8'hB1;
                    16'hECC6: data_out = 8'hB2;
                    16'hECC7: data_out = 8'hB3;
                    16'hECC8: data_out = 8'hB4;
                    16'hECC9: data_out = 8'hB5;
                    16'hECCA: data_out = 8'hB6;
                    16'hECCB: data_out = 8'hB7;
                    16'hECCC: data_out = 8'hB8;
                    16'hECCD: data_out = 8'hB9;
                    16'hECCE: data_out = 8'hBA;
                    16'hECCF: data_out = 8'hBB;
                    16'hECD0: data_out = 8'hBC;
                    16'hECD1: data_out = 8'hBD;
                    16'hECD2: data_out = 8'hBE;
                    16'hECD3: data_out = 8'hBF;
                    16'hECD4: data_out = 8'hC0;
                    16'hECD5: data_out = 8'hC1;
                    16'hECD6: data_out = 8'hC2;
                    16'hECD7: data_out = 8'hC3;
                    16'hECD8: data_out = 8'hC4;
                    16'hECD9: data_out = 8'hC5;
                    16'hECDA: data_out = 8'hC6;
                    16'hECDB: data_out = 8'hC7;
                    16'hECDC: data_out = 8'hC8;
                    16'hECDD: data_out = 8'hC9;
                    16'hECDE: data_out = 8'hCA;
                    16'hECDF: data_out = 8'hCB;
                    16'hECE0: data_out = 8'hCC;
                    16'hECE1: data_out = 8'hCD;
                    16'hECE2: data_out = 8'hCE;
                    16'hECE3: data_out = 8'hCF;
                    16'hECE4: data_out = 8'hD0;
                    16'hECE5: data_out = 8'hD1;
                    16'hECE6: data_out = 8'hD2;
                    16'hECE7: data_out = 8'hD3;
                    16'hECE8: data_out = 8'hD4;
                    16'hECE9: data_out = 8'hD5;
                    16'hECEA: data_out = 8'hD6;
                    16'hECEB: data_out = 8'hD7;
                    16'hECEC: data_out = 8'hD8;
                    16'hECED: data_out = 8'hD9;
                    16'hECEE: data_out = 8'hDA;
                    16'hECEF: data_out = 8'hDB;
                    16'hECF0: data_out = 8'hDC;
                    16'hECF1: data_out = 8'hDD;
                    16'hECF2: data_out = 8'hDE;
                    16'hECF3: data_out = 8'hDF;
                    16'hECF4: data_out = 8'hE0;
                    16'hECF5: data_out = 8'hE1;
                    16'hECF6: data_out = 8'hE2;
                    16'hECF7: data_out = 8'hE3;
                    16'hECF8: data_out = 8'hE4;
                    16'hECF9: data_out = 8'hE5;
                    16'hECFA: data_out = 8'hE6;
                    16'hECFB: data_out = 8'hE7;
                    16'hECFC: data_out = 8'hE8;
                    16'hECFD: data_out = 8'hE9;
                    16'hECFE: data_out = 8'hEA;
                    16'hECFF: data_out = 8'hEB;
                    16'hED00: data_out = 8'hED;
                    16'hED01: data_out = 8'hEC;
                    16'hED02: data_out = 8'hEB;
                    16'hED03: data_out = 8'hEA;
                    16'hED04: data_out = 8'hE9;
                    16'hED05: data_out = 8'hE8;
                    16'hED06: data_out = 8'hE7;
                    16'hED07: data_out = 8'hE6;
                    16'hED08: data_out = 8'hE5;
                    16'hED09: data_out = 8'hE4;
                    16'hED0A: data_out = 8'hE3;
                    16'hED0B: data_out = 8'hE2;
                    16'hED0C: data_out = 8'hE1;
                    16'hED0D: data_out = 8'hE0;
                    16'hED0E: data_out = 8'hDF;
                    16'hED0F: data_out = 8'hDE;
                    16'hED10: data_out = 8'hDD;
                    16'hED11: data_out = 8'hDC;
                    16'hED12: data_out = 8'hDB;
                    16'hED13: data_out = 8'hDA;
                    16'hED14: data_out = 8'hD9;
                    16'hED15: data_out = 8'hD8;
                    16'hED16: data_out = 8'hD7;
                    16'hED17: data_out = 8'hD6;
                    16'hED18: data_out = 8'hD5;
                    16'hED19: data_out = 8'hD4;
                    16'hED1A: data_out = 8'hD3;
                    16'hED1B: data_out = 8'hD2;
                    16'hED1C: data_out = 8'hD1;
                    16'hED1D: data_out = 8'hD0;
                    16'hED1E: data_out = 8'hCF;
                    16'hED1F: data_out = 8'hCE;
                    16'hED20: data_out = 8'hCD;
                    16'hED21: data_out = 8'hCC;
                    16'hED22: data_out = 8'hCB;
                    16'hED23: data_out = 8'hCA;
                    16'hED24: data_out = 8'hC9;
                    16'hED25: data_out = 8'hC8;
                    16'hED26: data_out = 8'hC7;
                    16'hED27: data_out = 8'hC6;
                    16'hED28: data_out = 8'hC5;
                    16'hED29: data_out = 8'hC4;
                    16'hED2A: data_out = 8'hC3;
                    16'hED2B: data_out = 8'hC2;
                    16'hED2C: data_out = 8'hC1;
                    16'hED2D: data_out = 8'hC0;
                    16'hED2E: data_out = 8'hBF;
                    16'hED2F: data_out = 8'hBE;
                    16'hED30: data_out = 8'hBD;
                    16'hED31: data_out = 8'hBC;
                    16'hED32: data_out = 8'hBB;
                    16'hED33: data_out = 8'hBA;
                    16'hED34: data_out = 8'hB9;
                    16'hED35: data_out = 8'hB8;
                    16'hED36: data_out = 8'hB7;
                    16'hED37: data_out = 8'hB6;
                    16'hED38: data_out = 8'hB5;
                    16'hED39: data_out = 8'hB4;
                    16'hED3A: data_out = 8'hB3;
                    16'hED3B: data_out = 8'hB2;
                    16'hED3C: data_out = 8'hB1;
                    16'hED3D: data_out = 8'hB0;
                    16'hED3E: data_out = 8'hAF;
                    16'hED3F: data_out = 8'hAE;
                    16'hED40: data_out = 8'hAD;
                    16'hED41: data_out = 8'hAC;
                    16'hED42: data_out = 8'hAB;
                    16'hED43: data_out = 8'hAA;
                    16'hED44: data_out = 8'hA9;
                    16'hED45: data_out = 8'hA8;
                    16'hED46: data_out = 8'hA7;
                    16'hED47: data_out = 8'hA6;
                    16'hED48: data_out = 8'hA5;
                    16'hED49: data_out = 8'hA4;
                    16'hED4A: data_out = 8'hA3;
                    16'hED4B: data_out = 8'hA2;
                    16'hED4C: data_out = 8'hA1;
                    16'hED4D: data_out = 8'hA0;
                    16'hED4E: data_out = 8'h9F;
                    16'hED4F: data_out = 8'h9E;
                    16'hED50: data_out = 8'h9D;
                    16'hED51: data_out = 8'h9C;
                    16'hED52: data_out = 8'h9B;
                    16'hED53: data_out = 8'h9A;
                    16'hED54: data_out = 8'h99;
                    16'hED55: data_out = 8'h98;
                    16'hED56: data_out = 8'h97;
                    16'hED57: data_out = 8'h96;
                    16'hED58: data_out = 8'h95;
                    16'hED59: data_out = 8'h94;
                    16'hED5A: data_out = 8'h93;
                    16'hED5B: data_out = 8'h92;
                    16'hED5C: data_out = 8'h91;
                    16'hED5D: data_out = 8'h90;
                    16'hED5E: data_out = 8'h8F;
                    16'hED5F: data_out = 8'h8E;
                    16'hED60: data_out = 8'h8D;
                    16'hED61: data_out = 8'h8C;
                    16'hED62: data_out = 8'h8B;
                    16'hED63: data_out = 8'h8A;
                    16'hED64: data_out = 8'h89;
                    16'hED65: data_out = 8'h88;
                    16'hED66: data_out = 8'h87;
                    16'hED67: data_out = 8'h86;
                    16'hED68: data_out = 8'h85;
                    16'hED69: data_out = 8'h84;
                    16'hED6A: data_out = 8'h83;
                    16'hED6B: data_out = 8'h82;
                    16'hED6C: data_out = 8'h81;
                    16'hED6D: data_out = 8'h0;
                    16'hED6E: data_out = 8'h1;
                    16'hED6F: data_out = 8'h2;
                    16'hED70: data_out = 8'h3;
                    16'hED71: data_out = 8'h4;
                    16'hED72: data_out = 8'h5;
                    16'hED73: data_out = 8'h6;
                    16'hED74: data_out = 8'h7;
                    16'hED75: data_out = 8'h8;
                    16'hED76: data_out = 8'h9;
                    16'hED77: data_out = 8'hA;
                    16'hED78: data_out = 8'hB;
                    16'hED79: data_out = 8'hC;
                    16'hED7A: data_out = 8'hD;
                    16'hED7B: data_out = 8'hE;
                    16'hED7C: data_out = 8'hF;
                    16'hED7D: data_out = 8'h10;
                    16'hED7E: data_out = 8'h11;
                    16'hED7F: data_out = 8'h12;
                    16'hED80: data_out = 8'hED;
                    16'hED81: data_out = 8'hEE;
                    16'hED82: data_out = 8'hEF;
                    16'hED83: data_out = 8'hF0;
                    16'hED84: data_out = 8'hF1;
                    16'hED85: data_out = 8'hF2;
                    16'hED86: data_out = 8'hF3;
                    16'hED87: data_out = 8'hF4;
                    16'hED88: data_out = 8'hF5;
                    16'hED89: data_out = 8'hF6;
                    16'hED8A: data_out = 8'hF7;
                    16'hED8B: data_out = 8'hF8;
                    16'hED8C: data_out = 8'hF9;
                    16'hED8D: data_out = 8'hFA;
                    16'hED8E: data_out = 8'hFB;
                    16'hED8F: data_out = 8'hFC;
                    16'hED90: data_out = 8'hFD;
                    16'hED91: data_out = 8'hFE;
                    16'hED92: data_out = 8'hFF;
                    16'hED93: data_out = 8'h80;
                    16'hED94: data_out = 8'h81;
                    16'hED95: data_out = 8'h82;
                    16'hED96: data_out = 8'h83;
                    16'hED97: data_out = 8'h84;
                    16'hED98: data_out = 8'h85;
                    16'hED99: data_out = 8'h86;
                    16'hED9A: data_out = 8'h87;
                    16'hED9B: data_out = 8'h88;
                    16'hED9C: data_out = 8'h89;
                    16'hED9D: data_out = 8'h8A;
                    16'hED9E: data_out = 8'h8B;
                    16'hED9F: data_out = 8'h8C;
                    16'hEDA0: data_out = 8'h8D;
                    16'hEDA1: data_out = 8'h8E;
                    16'hEDA2: data_out = 8'h8F;
                    16'hEDA3: data_out = 8'h90;
                    16'hEDA4: data_out = 8'h91;
                    16'hEDA5: data_out = 8'h92;
                    16'hEDA6: data_out = 8'h93;
                    16'hEDA7: data_out = 8'h94;
                    16'hEDA8: data_out = 8'h95;
                    16'hEDA9: data_out = 8'h96;
                    16'hEDAA: data_out = 8'h97;
                    16'hEDAB: data_out = 8'h98;
                    16'hEDAC: data_out = 8'h99;
                    16'hEDAD: data_out = 8'h9A;
                    16'hEDAE: data_out = 8'h9B;
                    16'hEDAF: data_out = 8'h9C;
                    16'hEDB0: data_out = 8'h9D;
                    16'hEDB1: data_out = 8'h9E;
                    16'hEDB2: data_out = 8'h9F;
                    16'hEDB3: data_out = 8'hA0;
                    16'hEDB4: data_out = 8'hA1;
                    16'hEDB5: data_out = 8'hA2;
                    16'hEDB6: data_out = 8'hA3;
                    16'hEDB7: data_out = 8'hA4;
                    16'hEDB8: data_out = 8'hA5;
                    16'hEDB9: data_out = 8'hA6;
                    16'hEDBA: data_out = 8'hA7;
                    16'hEDBB: data_out = 8'hA8;
                    16'hEDBC: data_out = 8'hA9;
                    16'hEDBD: data_out = 8'hAA;
                    16'hEDBE: data_out = 8'hAB;
                    16'hEDBF: data_out = 8'hAC;
                    16'hEDC0: data_out = 8'hAD;
                    16'hEDC1: data_out = 8'hAE;
                    16'hEDC2: data_out = 8'hAF;
                    16'hEDC3: data_out = 8'hB0;
                    16'hEDC4: data_out = 8'hB1;
                    16'hEDC5: data_out = 8'hB2;
                    16'hEDC6: data_out = 8'hB3;
                    16'hEDC7: data_out = 8'hB4;
                    16'hEDC8: data_out = 8'hB5;
                    16'hEDC9: data_out = 8'hB6;
                    16'hEDCA: data_out = 8'hB7;
                    16'hEDCB: data_out = 8'hB8;
                    16'hEDCC: data_out = 8'hB9;
                    16'hEDCD: data_out = 8'hBA;
                    16'hEDCE: data_out = 8'hBB;
                    16'hEDCF: data_out = 8'hBC;
                    16'hEDD0: data_out = 8'hBD;
                    16'hEDD1: data_out = 8'hBE;
                    16'hEDD2: data_out = 8'hBF;
                    16'hEDD3: data_out = 8'hC0;
                    16'hEDD4: data_out = 8'hC1;
                    16'hEDD5: data_out = 8'hC2;
                    16'hEDD6: data_out = 8'hC3;
                    16'hEDD7: data_out = 8'hC4;
                    16'hEDD8: data_out = 8'hC5;
                    16'hEDD9: data_out = 8'hC6;
                    16'hEDDA: data_out = 8'hC7;
                    16'hEDDB: data_out = 8'hC8;
                    16'hEDDC: data_out = 8'hC9;
                    16'hEDDD: data_out = 8'hCA;
                    16'hEDDE: data_out = 8'hCB;
                    16'hEDDF: data_out = 8'hCC;
                    16'hEDE0: data_out = 8'hCD;
                    16'hEDE1: data_out = 8'hCE;
                    16'hEDE2: data_out = 8'hCF;
                    16'hEDE3: data_out = 8'hD0;
                    16'hEDE4: data_out = 8'hD1;
                    16'hEDE5: data_out = 8'hD2;
                    16'hEDE6: data_out = 8'hD3;
                    16'hEDE7: data_out = 8'hD4;
                    16'hEDE8: data_out = 8'hD5;
                    16'hEDE9: data_out = 8'hD6;
                    16'hEDEA: data_out = 8'hD7;
                    16'hEDEB: data_out = 8'hD8;
                    16'hEDEC: data_out = 8'hD9;
                    16'hEDED: data_out = 8'hDA;
                    16'hEDEE: data_out = 8'hDB;
                    16'hEDEF: data_out = 8'hDC;
                    16'hEDF0: data_out = 8'hDD;
                    16'hEDF1: data_out = 8'hDE;
                    16'hEDF2: data_out = 8'hDF;
                    16'hEDF3: data_out = 8'hE0;
                    16'hEDF4: data_out = 8'hE1;
                    16'hEDF5: data_out = 8'hE2;
                    16'hEDF6: data_out = 8'hE3;
                    16'hEDF7: data_out = 8'hE4;
                    16'hEDF8: data_out = 8'hE5;
                    16'hEDF9: data_out = 8'hE6;
                    16'hEDFA: data_out = 8'hE7;
                    16'hEDFB: data_out = 8'hE8;
                    16'hEDFC: data_out = 8'hE9;
                    16'hEDFD: data_out = 8'hEA;
                    16'hEDFE: data_out = 8'hEB;
                    16'hEDFF: data_out = 8'hEC;
                    16'hEE00: data_out = 8'hEE;
                    16'hEE01: data_out = 8'hED;
                    16'hEE02: data_out = 8'hEC;
                    16'hEE03: data_out = 8'hEB;
                    16'hEE04: data_out = 8'hEA;
                    16'hEE05: data_out = 8'hE9;
                    16'hEE06: data_out = 8'hE8;
                    16'hEE07: data_out = 8'hE7;
                    16'hEE08: data_out = 8'hE6;
                    16'hEE09: data_out = 8'hE5;
                    16'hEE0A: data_out = 8'hE4;
                    16'hEE0B: data_out = 8'hE3;
                    16'hEE0C: data_out = 8'hE2;
                    16'hEE0D: data_out = 8'hE1;
                    16'hEE0E: data_out = 8'hE0;
                    16'hEE0F: data_out = 8'hDF;
                    16'hEE10: data_out = 8'hDE;
                    16'hEE11: data_out = 8'hDD;
                    16'hEE12: data_out = 8'hDC;
                    16'hEE13: data_out = 8'hDB;
                    16'hEE14: data_out = 8'hDA;
                    16'hEE15: data_out = 8'hD9;
                    16'hEE16: data_out = 8'hD8;
                    16'hEE17: data_out = 8'hD7;
                    16'hEE18: data_out = 8'hD6;
                    16'hEE19: data_out = 8'hD5;
                    16'hEE1A: data_out = 8'hD4;
                    16'hEE1B: data_out = 8'hD3;
                    16'hEE1C: data_out = 8'hD2;
                    16'hEE1D: data_out = 8'hD1;
                    16'hEE1E: data_out = 8'hD0;
                    16'hEE1F: data_out = 8'hCF;
                    16'hEE20: data_out = 8'hCE;
                    16'hEE21: data_out = 8'hCD;
                    16'hEE22: data_out = 8'hCC;
                    16'hEE23: data_out = 8'hCB;
                    16'hEE24: data_out = 8'hCA;
                    16'hEE25: data_out = 8'hC9;
                    16'hEE26: data_out = 8'hC8;
                    16'hEE27: data_out = 8'hC7;
                    16'hEE28: data_out = 8'hC6;
                    16'hEE29: data_out = 8'hC5;
                    16'hEE2A: data_out = 8'hC4;
                    16'hEE2B: data_out = 8'hC3;
                    16'hEE2C: data_out = 8'hC2;
                    16'hEE2D: data_out = 8'hC1;
                    16'hEE2E: data_out = 8'hC0;
                    16'hEE2F: data_out = 8'hBF;
                    16'hEE30: data_out = 8'hBE;
                    16'hEE31: data_out = 8'hBD;
                    16'hEE32: data_out = 8'hBC;
                    16'hEE33: data_out = 8'hBB;
                    16'hEE34: data_out = 8'hBA;
                    16'hEE35: data_out = 8'hB9;
                    16'hEE36: data_out = 8'hB8;
                    16'hEE37: data_out = 8'hB7;
                    16'hEE38: data_out = 8'hB6;
                    16'hEE39: data_out = 8'hB5;
                    16'hEE3A: data_out = 8'hB4;
                    16'hEE3B: data_out = 8'hB3;
                    16'hEE3C: data_out = 8'hB2;
                    16'hEE3D: data_out = 8'hB1;
                    16'hEE3E: data_out = 8'hB0;
                    16'hEE3F: data_out = 8'hAF;
                    16'hEE40: data_out = 8'hAE;
                    16'hEE41: data_out = 8'hAD;
                    16'hEE42: data_out = 8'hAC;
                    16'hEE43: data_out = 8'hAB;
                    16'hEE44: data_out = 8'hAA;
                    16'hEE45: data_out = 8'hA9;
                    16'hEE46: data_out = 8'hA8;
                    16'hEE47: data_out = 8'hA7;
                    16'hEE48: data_out = 8'hA6;
                    16'hEE49: data_out = 8'hA5;
                    16'hEE4A: data_out = 8'hA4;
                    16'hEE4B: data_out = 8'hA3;
                    16'hEE4C: data_out = 8'hA2;
                    16'hEE4D: data_out = 8'hA1;
                    16'hEE4E: data_out = 8'hA0;
                    16'hEE4F: data_out = 8'h9F;
                    16'hEE50: data_out = 8'h9E;
                    16'hEE51: data_out = 8'h9D;
                    16'hEE52: data_out = 8'h9C;
                    16'hEE53: data_out = 8'h9B;
                    16'hEE54: data_out = 8'h9A;
                    16'hEE55: data_out = 8'h99;
                    16'hEE56: data_out = 8'h98;
                    16'hEE57: data_out = 8'h97;
                    16'hEE58: data_out = 8'h96;
                    16'hEE59: data_out = 8'h95;
                    16'hEE5A: data_out = 8'h94;
                    16'hEE5B: data_out = 8'h93;
                    16'hEE5C: data_out = 8'h92;
                    16'hEE5D: data_out = 8'h91;
                    16'hEE5E: data_out = 8'h90;
                    16'hEE5F: data_out = 8'h8F;
                    16'hEE60: data_out = 8'h8E;
                    16'hEE61: data_out = 8'h8D;
                    16'hEE62: data_out = 8'h8C;
                    16'hEE63: data_out = 8'h8B;
                    16'hEE64: data_out = 8'h8A;
                    16'hEE65: data_out = 8'h89;
                    16'hEE66: data_out = 8'h88;
                    16'hEE67: data_out = 8'h87;
                    16'hEE68: data_out = 8'h86;
                    16'hEE69: data_out = 8'h85;
                    16'hEE6A: data_out = 8'h84;
                    16'hEE6B: data_out = 8'h83;
                    16'hEE6C: data_out = 8'h82;
                    16'hEE6D: data_out = 8'h81;
                    16'hEE6E: data_out = 8'h0;
                    16'hEE6F: data_out = 8'h1;
                    16'hEE70: data_out = 8'h2;
                    16'hEE71: data_out = 8'h3;
                    16'hEE72: data_out = 8'h4;
                    16'hEE73: data_out = 8'h5;
                    16'hEE74: data_out = 8'h6;
                    16'hEE75: data_out = 8'h7;
                    16'hEE76: data_out = 8'h8;
                    16'hEE77: data_out = 8'h9;
                    16'hEE78: data_out = 8'hA;
                    16'hEE79: data_out = 8'hB;
                    16'hEE7A: data_out = 8'hC;
                    16'hEE7B: data_out = 8'hD;
                    16'hEE7C: data_out = 8'hE;
                    16'hEE7D: data_out = 8'hF;
                    16'hEE7E: data_out = 8'h10;
                    16'hEE7F: data_out = 8'h11;
                    16'hEE80: data_out = 8'hEE;
                    16'hEE81: data_out = 8'hEF;
                    16'hEE82: data_out = 8'hF0;
                    16'hEE83: data_out = 8'hF1;
                    16'hEE84: data_out = 8'hF2;
                    16'hEE85: data_out = 8'hF3;
                    16'hEE86: data_out = 8'hF4;
                    16'hEE87: data_out = 8'hF5;
                    16'hEE88: data_out = 8'hF6;
                    16'hEE89: data_out = 8'hF7;
                    16'hEE8A: data_out = 8'hF8;
                    16'hEE8B: data_out = 8'hF9;
                    16'hEE8C: data_out = 8'hFA;
                    16'hEE8D: data_out = 8'hFB;
                    16'hEE8E: data_out = 8'hFC;
                    16'hEE8F: data_out = 8'hFD;
                    16'hEE90: data_out = 8'hFE;
                    16'hEE91: data_out = 8'hFF;
                    16'hEE92: data_out = 8'h80;
                    16'hEE93: data_out = 8'h81;
                    16'hEE94: data_out = 8'h82;
                    16'hEE95: data_out = 8'h83;
                    16'hEE96: data_out = 8'h84;
                    16'hEE97: data_out = 8'h85;
                    16'hEE98: data_out = 8'h86;
                    16'hEE99: data_out = 8'h87;
                    16'hEE9A: data_out = 8'h88;
                    16'hEE9B: data_out = 8'h89;
                    16'hEE9C: data_out = 8'h8A;
                    16'hEE9D: data_out = 8'h8B;
                    16'hEE9E: data_out = 8'h8C;
                    16'hEE9F: data_out = 8'h8D;
                    16'hEEA0: data_out = 8'h8E;
                    16'hEEA1: data_out = 8'h8F;
                    16'hEEA2: data_out = 8'h90;
                    16'hEEA3: data_out = 8'h91;
                    16'hEEA4: data_out = 8'h92;
                    16'hEEA5: data_out = 8'h93;
                    16'hEEA6: data_out = 8'h94;
                    16'hEEA7: data_out = 8'h95;
                    16'hEEA8: data_out = 8'h96;
                    16'hEEA9: data_out = 8'h97;
                    16'hEEAA: data_out = 8'h98;
                    16'hEEAB: data_out = 8'h99;
                    16'hEEAC: data_out = 8'h9A;
                    16'hEEAD: data_out = 8'h9B;
                    16'hEEAE: data_out = 8'h9C;
                    16'hEEAF: data_out = 8'h9D;
                    16'hEEB0: data_out = 8'h9E;
                    16'hEEB1: data_out = 8'h9F;
                    16'hEEB2: data_out = 8'hA0;
                    16'hEEB3: data_out = 8'hA1;
                    16'hEEB4: data_out = 8'hA2;
                    16'hEEB5: data_out = 8'hA3;
                    16'hEEB6: data_out = 8'hA4;
                    16'hEEB7: data_out = 8'hA5;
                    16'hEEB8: data_out = 8'hA6;
                    16'hEEB9: data_out = 8'hA7;
                    16'hEEBA: data_out = 8'hA8;
                    16'hEEBB: data_out = 8'hA9;
                    16'hEEBC: data_out = 8'hAA;
                    16'hEEBD: data_out = 8'hAB;
                    16'hEEBE: data_out = 8'hAC;
                    16'hEEBF: data_out = 8'hAD;
                    16'hEEC0: data_out = 8'hAE;
                    16'hEEC1: data_out = 8'hAF;
                    16'hEEC2: data_out = 8'hB0;
                    16'hEEC3: data_out = 8'hB1;
                    16'hEEC4: data_out = 8'hB2;
                    16'hEEC5: data_out = 8'hB3;
                    16'hEEC6: data_out = 8'hB4;
                    16'hEEC7: data_out = 8'hB5;
                    16'hEEC8: data_out = 8'hB6;
                    16'hEEC9: data_out = 8'hB7;
                    16'hEECA: data_out = 8'hB8;
                    16'hEECB: data_out = 8'hB9;
                    16'hEECC: data_out = 8'hBA;
                    16'hEECD: data_out = 8'hBB;
                    16'hEECE: data_out = 8'hBC;
                    16'hEECF: data_out = 8'hBD;
                    16'hEED0: data_out = 8'hBE;
                    16'hEED1: data_out = 8'hBF;
                    16'hEED2: data_out = 8'hC0;
                    16'hEED3: data_out = 8'hC1;
                    16'hEED4: data_out = 8'hC2;
                    16'hEED5: data_out = 8'hC3;
                    16'hEED6: data_out = 8'hC4;
                    16'hEED7: data_out = 8'hC5;
                    16'hEED8: data_out = 8'hC6;
                    16'hEED9: data_out = 8'hC7;
                    16'hEEDA: data_out = 8'hC8;
                    16'hEEDB: data_out = 8'hC9;
                    16'hEEDC: data_out = 8'hCA;
                    16'hEEDD: data_out = 8'hCB;
                    16'hEEDE: data_out = 8'hCC;
                    16'hEEDF: data_out = 8'hCD;
                    16'hEEE0: data_out = 8'hCE;
                    16'hEEE1: data_out = 8'hCF;
                    16'hEEE2: data_out = 8'hD0;
                    16'hEEE3: data_out = 8'hD1;
                    16'hEEE4: data_out = 8'hD2;
                    16'hEEE5: data_out = 8'hD3;
                    16'hEEE6: data_out = 8'hD4;
                    16'hEEE7: data_out = 8'hD5;
                    16'hEEE8: data_out = 8'hD6;
                    16'hEEE9: data_out = 8'hD7;
                    16'hEEEA: data_out = 8'hD8;
                    16'hEEEB: data_out = 8'hD9;
                    16'hEEEC: data_out = 8'hDA;
                    16'hEEED: data_out = 8'hDB;
                    16'hEEEE: data_out = 8'hDC;
                    16'hEEEF: data_out = 8'hDD;
                    16'hEEF0: data_out = 8'hDE;
                    16'hEEF1: data_out = 8'hDF;
                    16'hEEF2: data_out = 8'hE0;
                    16'hEEF3: data_out = 8'hE1;
                    16'hEEF4: data_out = 8'hE2;
                    16'hEEF5: data_out = 8'hE3;
                    16'hEEF6: data_out = 8'hE4;
                    16'hEEF7: data_out = 8'hE5;
                    16'hEEF8: data_out = 8'hE6;
                    16'hEEF9: data_out = 8'hE7;
                    16'hEEFA: data_out = 8'hE8;
                    16'hEEFB: data_out = 8'hE9;
                    16'hEEFC: data_out = 8'hEA;
                    16'hEEFD: data_out = 8'hEB;
                    16'hEEFE: data_out = 8'hEC;
                    16'hEEFF: data_out = 8'hED;
                    16'hEF00: data_out = 8'hEF;
                    16'hEF01: data_out = 8'hEE;
                    16'hEF02: data_out = 8'hED;
                    16'hEF03: data_out = 8'hEC;
                    16'hEF04: data_out = 8'hEB;
                    16'hEF05: data_out = 8'hEA;
                    16'hEF06: data_out = 8'hE9;
                    16'hEF07: data_out = 8'hE8;
                    16'hEF08: data_out = 8'hE7;
                    16'hEF09: data_out = 8'hE6;
                    16'hEF0A: data_out = 8'hE5;
                    16'hEF0B: data_out = 8'hE4;
                    16'hEF0C: data_out = 8'hE3;
                    16'hEF0D: data_out = 8'hE2;
                    16'hEF0E: data_out = 8'hE1;
                    16'hEF0F: data_out = 8'hE0;
                    16'hEF10: data_out = 8'hDF;
                    16'hEF11: data_out = 8'hDE;
                    16'hEF12: data_out = 8'hDD;
                    16'hEF13: data_out = 8'hDC;
                    16'hEF14: data_out = 8'hDB;
                    16'hEF15: data_out = 8'hDA;
                    16'hEF16: data_out = 8'hD9;
                    16'hEF17: data_out = 8'hD8;
                    16'hEF18: data_out = 8'hD7;
                    16'hEF19: data_out = 8'hD6;
                    16'hEF1A: data_out = 8'hD5;
                    16'hEF1B: data_out = 8'hD4;
                    16'hEF1C: data_out = 8'hD3;
                    16'hEF1D: data_out = 8'hD2;
                    16'hEF1E: data_out = 8'hD1;
                    16'hEF1F: data_out = 8'hD0;
                    16'hEF20: data_out = 8'hCF;
                    16'hEF21: data_out = 8'hCE;
                    16'hEF22: data_out = 8'hCD;
                    16'hEF23: data_out = 8'hCC;
                    16'hEF24: data_out = 8'hCB;
                    16'hEF25: data_out = 8'hCA;
                    16'hEF26: data_out = 8'hC9;
                    16'hEF27: data_out = 8'hC8;
                    16'hEF28: data_out = 8'hC7;
                    16'hEF29: data_out = 8'hC6;
                    16'hEF2A: data_out = 8'hC5;
                    16'hEF2B: data_out = 8'hC4;
                    16'hEF2C: data_out = 8'hC3;
                    16'hEF2D: data_out = 8'hC2;
                    16'hEF2E: data_out = 8'hC1;
                    16'hEF2F: data_out = 8'hC0;
                    16'hEF30: data_out = 8'hBF;
                    16'hEF31: data_out = 8'hBE;
                    16'hEF32: data_out = 8'hBD;
                    16'hEF33: data_out = 8'hBC;
                    16'hEF34: data_out = 8'hBB;
                    16'hEF35: data_out = 8'hBA;
                    16'hEF36: data_out = 8'hB9;
                    16'hEF37: data_out = 8'hB8;
                    16'hEF38: data_out = 8'hB7;
                    16'hEF39: data_out = 8'hB6;
                    16'hEF3A: data_out = 8'hB5;
                    16'hEF3B: data_out = 8'hB4;
                    16'hEF3C: data_out = 8'hB3;
                    16'hEF3D: data_out = 8'hB2;
                    16'hEF3E: data_out = 8'hB1;
                    16'hEF3F: data_out = 8'hB0;
                    16'hEF40: data_out = 8'hAF;
                    16'hEF41: data_out = 8'hAE;
                    16'hEF42: data_out = 8'hAD;
                    16'hEF43: data_out = 8'hAC;
                    16'hEF44: data_out = 8'hAB;
                    16'hEF45: data_out = 8'hAA;
                    16'hEF46: data_out = 8'hA9;
                    16'hEF47: data_out = 8'hA8;
                    16'hEF48: data_out = 8'hA7;
                    16'hEF49: data_out = 8'hA6;
                    16'hEF4A: data_out = 8'hA5;
                    16'hEF4B: data_out = 8'hA4;
                    16'hEF4C: data_out = 8'hA3;
                    16'hEF4D: data_out = 8'hA2;
                    16'hEF4E: data_out = 8'hA1;
                    16'hEF4F: data_out = 8'hA0;
                    16'hEF50: data_out = 8'h9F;
                    16'hEF51: data_out = 8'h9E;
                    16'hEF52: data_out = 8'h9D;
                    16'hEF53: data_out = 8'h9C;
                    16'hEF54: data_out = 8'h9B;
                    16'hEF55: data_out = 8'h9A;
                    16'hEF56: data_out = 8'h99;
                    16'hEF57: data_out = 8'h98;
                    16'hEF58: data_out = 8'h97;
                    16'hEF59: data_out = 8'h96;
                    16'hEF5A: data_out = 8'h95;
                    16'hEF5B: data_out = 8'h94;
                    16'hEF5C: data_out = 8'h93;
                    16'hEF5D: data_out = 8'h92;
                    16'hEF5E: data_out = 8'h91;
                    16'hEF5F: data_out = 8'h90;
                    16'hEF60: data_out = 8'h8F;
                    16'hEF61: data_out = 8'h8E;
                    16'hEF62: data_out = 8'h8D;
                    16'hEF63: data_out = 8'h8C;
                    16'hEF64: data_out = 8'h8B;
                    16'hEF65: data_out = 8'h8A;
                    16'hEF66: data_out = 8'h89;
                    16'hEF67: data_out = 8'h88;
                    16'hEF68: data_out = 8'h87;
                    16'hEF69: data_out = 8'h86;
                    16'hEF6A: data_out = 8'h85;
                    16'hEF6B: data_out = 8'h84;
                    16'hEF6C: data_out = 8'h83;
                    16'hEF6D: data_out = 8'h82;
                    16'hEF6E: data_out = 8'h81;
                    16'hEF6F: data_out = 8'h0;
                    16'hEF70: data_out = 8'h1;
                    16'hEF71: data_out = 8'h2;
                    16'hEF72: data_out = 8'h3;
                    16'hEF73: data_out = 8'h4;
                    16'hEF74: data_out = 8'h5;
                    16'hEF75: data_out = 8'h6;
                    16'hEF76: data_out = 8'h7;
                    16'hEF77: data_out = 8'h8;
                    16'hEF78: data_out = 8'h9;
                    16'hEF79: data_out = 8'hA;
                    16'hEF7A: data_out = 8'hB;
                    16'hEF7B: data_out = 8'hC;
                    16'hEF7C: data_out = 8'hD;
                    16'hEF7D: data_out = 8'hE;
                    16'hEF7E: data_out = 8'hF;
                    16'hEF7F: data_out = 8'h10;
                    16'hEF80: data_out = 8'hEF;
                    16'hEF81: data_out = 8'hF0;
                    16'hEF82: data_out = 8'hF1;
                    16'hEF83: data_out = 8'hF2;
                    16'hEF84: data_out = 8'hF3;
                    16'hEF85: data_out = 8'hF4;
                    16'hEF86: data_out = 8'hF5;
                    16'hEF87: data_out = 8'hF6;
                    16'hEF88: data_out = 8'hF7;
                    16'hEF89: data_out = 8'hF8;
                    16'hEF8A: data_out = 8'hF9;
                    16'hEF8B: data_out = 8'hFA;
                    16'hEF8C: data_out = 8'hFB;
                    16'hEF8D: data_out = 8'hFC;
                    16'hEF8E: data_out = 8'hFD;
                    16'hEF8F: data_out = 8'hFE;
                    16'hEF90: data_out = 8'hFF;
                    16'hEF91: data_out = 8'h80;
                    16'hEF92: data_out = 8'h81;
                    16'hEF93: data_out = 8'h82;
                    16'hEF94: data_out = 8'h83;
                    16'hEF95: data_out = 8'h84;
                    16'hEF96: data_out = 8'h85;
                    16'hEF97: data_out = 8'h86;
                    16'hEF98: data_out = 8'h87;
                    16'hEF99: data_out = 8'h88;
                    16'hEF9A: data_out = 8'h89;
                    16'hEF9B: data_out = 8'h8A;
                    16'hEF9C: data_out = 8'h8B;
                    16'hEF9D: data_out = 8'h8C;
                    16'hEF9E: data_out = 8'h8D;
                    16'hEF9F: data_out = 8'h8E;
                    16'hEFA0: data_out = 8'h8F;
                    16'hEFA1: data_out = 8'h90;
                    16'hEFA2: data_out = 8'h91;
                    16'hEFA3: data_out = 8'h92;
                    16'hEFA4: data_out = 8'h93;
                    16'hEFA5: data_out = 8'h94;
                    16'hEFA6: data_out = 8'h95;
                    16'hEFA7: data_out = 8'h96;
                    16'hEFA8: data_out = 8'h97;
                    16'hEFA9: data_out = 8'h98;
                    16'hEFAA: data_out = 8'h99;
                    16'hEFAB: data_out = 8'h9A;
                    16'hEFAC: data_out = 8'h9B;
                    16'hEFAD: data_out = 8'h9C;
                    16'hEFAE: data_out = 8'h9D;
                    16'hEFAF: data_out = 8'h9E;
                    16'hEFB0: data_out = 8'h9F;
                    16'hEFB1: data_out = 8'hA0;
                    16'hEFB2: data_out = 8'hA1;
                    16'hEFB3: data_out = 8'hA2;
                    16'hEFB4: data_out = 8'hA3;
                    16'hEFB5: data_out = 8'hA4;
                    16'hEFB6: data_out = 8'hA5;
                    16'hEFB7: data_out = 8'hA6;
                    16'hEFB8: data_out = 8'hA7;
                    16'hEFB9: data_out = 8'hA8;
                    16'hEFBA: data_out = 8'hA9;
                    16'hEFBB: data_out = 8'hAA;
                    16'hEFBC: data_out = 8'hAB;
                    16'hEFBD: data_out = 8'hAC;
                    16'hEFBE: data_out = 8'hAD;
                    16'hEFBF: data_out = 8'hAE;
                    16'hEFC0: data_out = 8'hAF;
                    16'hEFC1: data_out = 8'hB0;
                    16'hEFC2: data_out = 8'hB1;
                    16'hEFC3: data_out = 8'hB2;
                    16'hEFC4: data_out = 8'hB3;
                    16'hEFC5: data_out = 8'hB4;
                    16'hEFC6: data_out = 8'hB5;
                    16'hEFC7: data_out = 8'hB6;
                    16'hEFC8: data_out = 8'hB7;
                    16'hEFC9: data_out = 8'hB8;
                    16'hEFCA: data_out = 8'hB9;
                    16'hEFCB: data_out = 8'hBA;
                    16'hEFCC: data_out = 8'hBB;
                    16'hEFCD: data_out = 8'hBC;
                    16'hEFCE: data_out = 8'hBD;
                    16'hEFCF: data_out = 8'hBE;
                    16'hEFD0: data_out = 8'hBF;
                    16'hEFD1: data_out = 8'hC0;
                    16'hEFD2: data_out = 8'hC1;
                    16'hEFD3: data_out = 8'hC2;
                    16'hEFD4: data_out = 8'hC3;
                    16'hEFD5: data_out = 8'hC4;
                    16'hEFD6: data_out = 8'hC5;
                    16'hEFD7: data_out = 8'hC6;
                    16'hEFD8: data_out = 8'hC7;
                    16'hEFD9: data_out = 8'hC8;
                    16'hEFDA: data_out = 8'hC9;
                    16'hEFDB: data_out = 8'hCA;
                    16'hEFDC: data_out = 8'hCB;
                    16'hEFDD: data_out = 8'hCC;
                    16'hEFDE: data_out = 8'hCD;
                    16'hEFDF: data_out = 8'hCE;
                    16'hEFE0: data_out = 8'hCF;
                    16'hEFE1: data_out = 8'hD0;
                    16'hEFE2: data_out = 8'hD1;
                    16'hEFE3: data_out = 8'hD2;
                    16'hEFE4: data_out = 8'hD3;
                    16'hEFE5: data_out = 8'hD4;
                    16'hEFE6: data_out = 8'hD5;
                    16'hEFE7: data_out = 8'hD6;
                    16'hEFE8: data_out = 8'hD7;
                    16'hEFE9: data_out = 8'hD8;
                    16'hEFEA: data_out = 8'hD9;
                    16'hEFEB: data_out = 8'hDA;
                    16'hEFEC: data_out = 8'hDB;
                    16'hEFED: data_out = 8'hDC;
                    16'hEFEE: data_out = 8'hDD;
                    16'hEFEF: data_out = 8'hDE;
                    16'hEFF0: data_out = 8'hDF;
                    16'hEFF1: data_out = 8'hE0;
                    16'hEFF2: data_out = 8'hE1;
                    16'hEFF3: data_out = 8'hE2;
                    16'hEFF4: data_out = 8'hE3;
                    16'hEFF5: data_out = 8'hE4;
                    16'hEFF6: data_out = 8'hE5;
                    16'hEFF7: data_out = 8'hE6;
                    16'hEFF8: data_out = 8'hE7;
                    16'hEFF9: data_out = 8'hE8;
                    16'hEFFA: data_out = 8'hE9;
                    16'hEFFB: data_out = 8'hEA;
                    16'hEFFC: data_out = 8'hEB;
                    16'hEFFD: data_out = 8'hEC;
                    16'hEFFE: data_out = 8'hED;
                    16'hEFFF: data_out = 8'hEE;
                    16'hF000: data_out = 8'hF0;
                    16'hF001: data_out = 8'hEF;
                    16'hF002: data_out = 8'hEE;
                    16'hF003: data_out = 8'hED;
                    16'hF004: data_out = 8'hEC;
                    16'hF005: data_out = 8'hEB;
                    16'hF006: data_out = 8'hEA;
                    16'hF007: data_out = 8'hE9;
                    16'hF008: data_out = 8'hE8;
                    16'hF009: data_out = 8'hE7;
                    16'hF00A: data_out = 8'hE6;
                    16'hF00B: data_out = 8'hE5;
                    16'hF00C: data_out = 8'hE4;
                    16'hF00D: data_out = 8'hE3;
                    16'hF00E: data_out = 8'hE2;
                    16'hF00F: data_out = 8'hE1;
                    16'hF010: data_out = 8'hE0;
                    16'hF011: data_out = 8'hDF;
                    16'hF012: data_out = 8'hDE;
                    16'hF013: data_out = 8'hDD;
                    16'hF014: data_out = 8'hDC;
                    16'hF015: data_out = 8'hDB;
                    16'hF016: data_out = 8'hDA;
                    16'hF017: data_out = 8'hD9;
                    16'hF018: data_out = 8'hD8;
                    16'hF019: data_out = 8'hD7;
                    16'hF01A: data_out = 8'hD6;
                    16'hF01B: data_out = 8'hD5;
                    16'hF01C: data_out = 8'hD4;
                    16'hF01D: data_out = 8'hD3;
                    16'hF01E: data_out = 8'hD2;
                    16'hF01F: data_out = 8'hD1;
                    16'hF020: data_out = 8'hD0;
                    16'hF021: data_out = 8'hCF;
                    16'hF022: data_out = 8'hCE;
                    16'hF023: data_out = 8'hCD;
                    16'hF024: data_out = 8'hCC;
                    16'hF025: data_out = 8'hCB;
                    16'hF026: data_out = 8'hCA;
                    16'hF027: data_out = 8'hC9;
                    16'hF028: data_out = 8'hC8;
                    16'hF029: data_out = 8'hC7;
                    16'hF02A: data_out = 8'hC6;
                    16'hF02B: data_out = 8'hC5;
                    16'hF02C: data_out = 8'hC4;
                    16'hF02D: data_out = 8'hC3;
                    16'hF02E: data_out = 8'hC2;
                    16'hF02F: data_out = 8'hC1;
                    16'hF030: data_out = 8'hC0;
                    16'hF031: data_out = 8'hBF;
                    16'hF032: data_out = 8'hBE;
                    16'hF033: data_out = 8'hBD;
                    16'hF034: data_out = 8'hBC;
                    16'hF035: data_out = 8'hBB;
                    16'hF036: data_out = 8'hBA;
                    16'hF037: data_out = 8'hB9;
                    16'hF038: data_out = 8'hB8;
                    16'hF039: data_out = 8'hB7;
                    16'hF03A: data_out = 8'hB6;
                    16'hF03B: data_out = 8'hB5;
                    16'hF03C: data_out = 8'hB4;
                    16'hF03D: data_out = 8'hB3;
                    16'hF03E: data_out = 8'hB2;
                    16'hF03F: data_out = 8'hB1;
                    16'hF040: data_out = 8'hB0;
                    16'hF041: data_out = 8'hAF;
                    16'hF042: data_out = 8'hAE;
                    16'hF043: data_out = 8'hAD;
                    16'hF044: data_out = 8'hAC;
                    16'hF045: data_out = 8'hAB;
                    16'hF046: data_out = 8'hAA;
                    16'hF047: data_out = 8'hA9;
                    16'hF048: data_out = 8'hA8;
                    16'hF049: data_out = 8'hA7;
                    16'hF04A: data_out = 8'hA6;
                    16'hF04B: data_out = 8'hA5;
                    16'hF04C: data_out = 8'hA4;
                    16'hF04D: data_out = 8'hA3;
                    16'hF04E: data_out = 8'hA2;
                    16'hF04F: data_out = 8'hA1;
                    16'hF050: data_out = 8'hA0;
                    16'hF051: data_out = 8'h9F;
                    16'hF052: data_out = 8'h9E;
                    16'hF053: data_out = 8'h9D;
                    16'hF054: data_out = 8'h9C;
                    16'hF055: data_out = 8'h9B;
                    16'hF056: data_out = 8'h9A;
                    16'hF057: data_out = 8'h99;
                    16'hF058: data_out = 8'h98;
                    16'hF059: data_out = 8'h97;
                    16'hF05A: data_out = 8'h96;
                    16'hF05B: data_out = 8'h95;
                    16'hF05C: data_out = 8'h94;
                    16'hF05D: data_out = 8'h93;
                    16'hF05E: data_out = 8'h92;
                    16'hF05F: data_out = 8'h91;
                    16'hF060: data_out = 8'h90;
                    16'hF061: data_out = 8'h8F;
                    16'hF062: data_out = 8'h8E;
                    16'hF063: data_out = 8'h8D;
                    16'hF064: data_out = 8'h8C;
                    16'hF065: data_out = 8'h8B;
                    16'hF066: data_out = 8'h8A;
                    16'hF067: data_out = 8'h89;
                    16'hF068: data_out = 8'h88;
                    16'hF069: data_out = 8'h87;
                    16'hF06A: data_out = 8'h86;
                    16'hF06B: data_out = 8'h85;
                    16'hF06C: data_out = 8'h84;
                    16'hF06D: data_out = 8'h83;
                    16'hF06E: data_out = 8'h82;
                    16'hF06F: data_out = 8'h81;
                    16'hF070: data_out = 8'h0;
                    16'hF071: data_out = 8'h1;
                    16'hF072: data_out = 8'h2;
                    16'hF073: data_out = 8'h3;
                    16'hF074: data_out = 8'h4;
                    16'hF075: data_out = 8'h5;
                    16'hF076: data_out = 8'h6;
                    16'hF077: data_out = 8'h7;
                    16'hF078: data_out = 8'h8;
                    16'hF079: data_out = 8'h9;
                    16'hF07A: data_out = 8'hA;
                    16'hF07B: data_out = 8'hB;
                    16'hF07C: data_out = 8'hC;
                    16'hF07D: data_out = 8'hD;
                    16'hF07E: data_out = 8'hE;
                    16'hF07F: data_out = 8'hF;
                    16'hF080: data_out = 8'hF0;
                    16'hF081: data_out = 8'hF1;
                    16'hF082: data_out = 8'hF2;
                    16'hF083: data_out = 8'hF3;
                    16'hF084: data_out = 8'hF4;
                    16'hF085: data_out = 8'hF5;
                    16'hF086: data_out = 8'hF6;
                    16'hF087: data_out = 8'hF7;
                    16'hF088: data_out = 8'hF8;
                    16'hF089: data_out = 8'hF9;
                    16'hF08A: data_out = 8'hFA;
                    16'hF08B: data_out = 8'hFB;
                    16'hF08C: data_out = 8'hFC;
                    16'hF08D: data_out = 8'hFD;
                    16'hF08E: data_out = 8'hFE;
                    16'hF08F: data_out = 8'hFF;
                    16'hF090: data_out = 8'h80;
                    16'hF091: data_out = 8'h81;
                    16'hF092: data_out = 8'h82;
                    16'hF093: data_out = 8'h83;
                    16'hF094: data_out = 8'h84;
                    16'hF095: data_out = 8'h85;
                    16'hF096: data_out = 8'h86;
                    16'hF097: data_out = 8'h87;
                    16'hF098: data_out = 8'h88;
                    16'hF099: data_out = 8'h89;
                    16'hF09A: data_out = 8'h8A;
                    16'hF09B: data_out = 8'h8B;
                    16'hF09C: data_out = 8'h8C;
                    16'hF09D: data_out = 8'h8D;
                    16'hF09E: data_out = 8'h8E;
                    16'hF09F: data_out = 8'h8F;
                    16'hF0A0: data_out = 8'h90;
                    16'hF0A1: data_out = 8'h91;
                    16'hF0A2: data_out = 8'h92;
                    16'hF0A3: data_out = 8'h93;
                    16'hF0A4: data_out = 8'h94;
                    16'hF0A5: data_out = 8'h95;
                    16'hF0A6: data_out = 8'h96;
                    16'hF0A7: data_out = 8'h97;
                    16'hF0A8: data_out = 8'h98;
                    16'hF0A9: data_out = 8'h99;
                    16'hF0AA: data_out = 8'h9A;
                    16'hF0AB: data_out = 8'h9B;
                    16'hF0AC: data_out = 8'h9C;
                    16'hF0AD: data_out = 8'h9D;
                    16'hF0AE: data_out = 8'h9E;
                    16'hF0AF: data_out = 8'h9F;
                    16'hF0B0: data_out = 8'hA0;
                    16'hF0B1: data_out = 8'hA1;
                    16'hF0B2: data_out = 8'hA2;
                    16'hF0B3: data_out = 8'hA3;
                    16'hF0B4: data_out = 8'hA4;
                    16'hF0B5: data_out = 8'hA5;
                    16'hF0B6: data_out = 8'hA6;
                    16'hF0B7: data_out = 8'hA7;
                    16'hF0B8: data_out = 8'hA8;
                    16'hF0B9: data_out = 8'hA9;
                    16'hF0BA: data_out = 8'hAA;
                    16'hF0BB: data_out = 8'hAB;
                    16'hF0BC: data_out = 8'hAC;
                    16'hF0BD: data_out = 8'hAD;
                    16'hF0BE: data_out = 8'hAE;
                    16'hF0BF: data_out = 8'hAF;
                    16'hF0C0: data_out = 8'hB0;
                    16'hF0C1: data_out = 8'hB1;
                    16'hF0C2: data_out = 8'hB2;
                    16'hF0C3: data_out = 8'hB3;
                    16'hF0C4: data_out = 8'hB4;
                    16'hF0C5: data_out = 8'hB5;
                    16'hF0C6: data_out = 8'hB6;
                    16'hF0C7: data_out = 8'hB7;
                    16'hF0C8: data_out = 8'hB8;
                    16'hF0C9: data_out = 8'hB9;
                    16'hF0CA: data_out = 8'hBA;
                    16'hF0CB: data_out = 8'hBB;
                    16'hF0CC: data_out = 8'hBC;
                    16'hF0CD: data_out = 8'hBD;
                    16'hF0CE: data_out = 8'hBE;
                    16'hF0CF: data_out = 8'hBF;
                    16'hF0D0: data_out = 8'hC0;
                    16'hF0D1: data_out = 8'hC1;
                    16'hF0D2: data_out = 8'hC2;
                    16'hF0D3: data_out = 8'hC3;
                    16'hF0D4: data_out = 8'hC4;
                    16'hF0D5: data_out = 8'hC5;
                    16'hF0D6: data_out = 8'hC6;
                    16'hF0D7: data_out = 8'hC7;
                    16'hF0D8: data_out = 8'hC8;
                    16'hF0D9: data_out = 8'hC9;
                    16'hF0DA: data_out = 8'hCA;
                    16'hF0DB: data_out = 8'hCB;
                    16'hF0DC: data_out = 8'hCC;
                    16'hF0DD: data_out = 8'hCD;
                    16'hF0DE: data_out = 8'hCE;
                    16'hF0DF: data_out = 8'hCF;
                    16'hF0E0: data_out = 8'hD0;
                    16'hF0E1: data_out = 8'hD1;
                    16'hF0E2: data_out = 8'hD2;
                    16'hF0E3: data_out = 8'hD3;
                    16'hF0E4: data_out = 8'hD4;
                    16'hF0E5: data_out = 8'hD5;
                    16'hF0E6: data_out = 8'hD6;
                    16'hF0E7: data_out = 8'hD7;
                    16'hF0E8: data_out = 8'hD8;
                    16'hF0E9: data_out = 8'hD9;
                    16'hF0EA: data_out = 8'hDA;
                    16'hF0EB: data_out = 8'hDB;
                    16'hF0EC: data_out = 8'hDC;
                    16'hF0ED: data_out = 8'hDD;
                    16'hF0EE: data_out = 8'hDE;
                    16'hF0EF: data_out = 8'hDF;
                    16'hF0F0: data_out = 8'hE0;
                    16'hF0F1: data_out = 8'hE1;
                    16'hF0F2: data_out = 8'hE2;
                    16'hF0F3: data_out = 8'hE3;
                    16'hF0F4: data_out = 8'hE4;
                    16'hF0F5: data_out = 8'hE5;
                    16'hF0F6: data_out = 8'hE6;
                    16'hF0F7: data_out = 8'hE7;
                    16'hF0F8: data_out = 8'hE8;
                    16'hF0F9: data_out = 8'hE9;
                    16'hF0FA: data_out = 8'hEA;
                    16'hF0FB: data_out = 8'hEB;
                    16'hF0FC: data_out = 8'hEC;
                    16'hF0FD: data_out = 8'hED;
                    16'hF0FE: data_out = 8'hEE;
                    16'hF0FF: data_out = 8'hEF;
                    16'hF100: data_out = 8'hF1;
                    16'hF101: data_out = 8'hF0;
                    16'hF102: data_out = 8'hEF;
                    16'hF103: data_out = 8'hEE;
                    16'hF104: data_out = 8'hED;
                    16'hF105: data_out = 8'hEC;
                    16'hF106: data_out = 8'hEB;
                    16'hF107: data_out = 8'hEA;
                    16'hF108: data_out = 8'hE9;
                    16'hF109: data_out = 8'hE8;
                    16'hF10A: data_out = 8'hE7;
                    16'hF10B: data_out = 8'hE6;
                    16'hF10C: data_out = 8'hE5;
                    16'hF10D: data_out = 8'hE4;
                    16'hF10E: data_out = 8'hE3;
                    16'hF10F: data_out = 8'hE2;
                    16'hF110: data_out = 8'hE1;
                    16'hF111: data_out = 8'hE0;
                    16'hF112: data_out = 8'hDF;
                    16'hF113: data_out = 8'hDE;
                    16'hF114: data_out = 8'hDD;
                    16'hF115: data_out = 8'hDC;
                    16'hF116: data_out = 8'hDB;
                    16'hF117: data_out = 8'hDA;
                    16'hF118: data_out = 8'hD9;
                    16'hF119: data_out = 8'hD8;
                    16'hF11A: data_out = 8'hD7;
                    16'hF11B: data_out = 8'hD6;
                    16'hF11C: data_out = 8'hD5;
                    16'hF11D: data_out = 8'hD4;
                    16'hF11E: data_out = 8'hD3;
                    16'hF11F: data_out = 8'hD2;
                    16'hF120: data_out = 8'hD1;
                    16'hF121: data_out = 8'hD0;
                    16'hF122: data_out = 8'hCF;
                    16'hF123: data_out = 8'hCE;
                    16'hF124: data_out = 8'hCD;
                    16'hF125: data_out = 8'hCC;
                    16'hF126: data_out = 8'hCB;
                    16'hF127: data_out = 8'hCA;
                    16'hF128: data_out = 8'hC9;
                    16'hF129: data_out = 8'hC8;
                    16'hF12A: data_out = 8'hC7;
                    16'hF12B: data_out = 8'hC6;
                    16'hF12C: data_out = 8'hC5;
                    16'hF12D: data_out = 8'hC4;
                    16'hF12E: data_out = 8'hC3;
                    16'hF12F: data_out = 8'hC2;
                    16'hF130: data_out = 8'hC1;
                    16'hF131: data_out = 8'hC0;
                    16'hF132: data_out = 8'hBF;
                    16'hF133: data_out = 8'hBE;
                    16'hF134: data_out = 8'hBD;
                    16'hF135: data_out = 8'hBC;
                    16'hF136: data_out = 8'hBB;
                    16'hF137: data_out = 8'hBA;
                    16'hF138: data_out = 8'hB9;
                    16'hF139: data_out = 8'hB8;
                    16'hF13A: data_out = 8'hB7;
                    16'hF13B: data_out = 8'hB6;
                    16'hF13C: data_out = 8'hB5;
                    16'hF13D: data_out = 8'hB4;
                    16'hF13E: data_out = 8'hB3;
                    16'hF13F: data_out = 8'hB2;
                    16'hF140: data_out = 8'hB1;
                    16'hF141: data_out = 8'hB0;
                    16'hF142: data_out = 8'hAF;
                    16'hF143: data_out = 8'hAE;
                    16'hF144: data_out = 8'hAD;
                    16'hF145: data_out = 8'hAC;
                    16'hF146: data_out = 8'hAB;
                    16'hF147: data_out = 8'hAA;
                    16'hF148: data_out = 8'hA9;
                    16'hF149: data_out = 8'hA8;
                    16'hF14A: data_out = 8'hA7;
                    16'hF14B: data_out = 8'hA6;
                    16'hF14C: data_out = 8'hA5;
                    16'hF14D: data_out = 8'hA4;
                    16'hF14E: data_out = 8'hA3;
                    16'hF14F: data_out = 8'hA2;
                    16'hF150: data_out = 8'hA1;
                    16'hF151: data_out = 8'hA0;
                    16'hF152: data_out = 8'h9F;
                    16'hF153: data_out = 8'h9E;
                    16'hF154: data_out = 8'h9D;
                    16'hF155: data_out = 8'h9C;
                    16'hF156: data_out = 8'h9B;
                    16'hF157: data_out = 8'h9A;
                    16'hF158: data_out = 8'h99;
                    16'hF159: data_out = 8'h98;
                    16'hF15A: data_out = 8'h97;
                    16'hF15B: data_out = 8'h96;
                    16'hF15C: data_out = 8'h95;
                    16'hF15D: data_out = 8'h94;
                    16'hF15E: data_out = 8'h93;
                    16'hF15F: data_out = 8'h92;
                    16'hF160: data_out = 8'h91;
                    16'hF161: data_out = 8'h90;
                    16'hF162: data_out = 8'h8F;
                    16'hF163: data_out = 8'h8E;
                    16'hF164: data_out = 8'h8D;
                    16'hF165: data_out = 8'h8C;
                    16'hF166: data_out = 8'h8B;
                    16'hF167: data_out = 8'h8A;
                    16'hF168: data_out = 8'h89;
                    16'hF169: data_out = 8'h88;
                    16'hF16A: data_out = 8'h87;
                    16'hF16B: data_out = 8'h86;
                    16'hF16C: data_out = 8'h85;
                    16'hF16D: data_out = 8'h84;
                    16'hF16E: data_out = 8'h83;
                    16'hF16F: data_out = 8'h82;
                    16'hF170: data_out = 8'h81;
                    16'hF171: data_out = 8'h0;
                    16'hF172: data_out = 8'h1;
                    16'hF173: data_out = 8'h2;
                    16'hF174: data_out = 8'h3;
                    16'hF175: data_out = 8'h4;
                    16'hF176: data_out = 8'h5;
                    16'hF177: data_out = 8'h6;
                    16'hF178: data_out = 8'h7;
                    16'hF179: data_out = 8'h8;
                    16'hF17A: data_out = 8'h9;
                    16'hF17B: data_out = 8'hA;
                    16'hF17C: data_out = 8'hB;
                    16'hF17D: data_out = 8'hC;
                    16'hF17E: data_out = 8'hD;
                    16'hF17F: data_out = 8'hE;
                    16'hF180: data_out = 8'hF1;
                    16'hF181: data_out = 8'hF2;
                    16'hF182: data_out = 8'hF3;
                    16'hF183: data_out = 8'hF4;
                    16'hF184: data_out = 8'hF5;
                    16'hF185: data_out = 8'hF6;
                    16'hF186: data_out = 8'hF7;
                    16'hF187: data_out = 8'hF8;
                    16'hF188: data_out = 8'hF9;
                    16'hF189: data_out = 8'hFA;
                    16'hF18A: data_out = 8'hFB;
                    16'hF18B: data_out = 8'hFC;
                    16'hF18C: data_out = 8'hFD;
                    16'hF18D: data_out = 8'hFE;
                    16'hF18E: data_out = 8'hFF;
                    16'hF18F: data_out = 8'h80;
                    16'hF190: data_out = 8'h81;
                    16'hF191: data_out = 8'h82;
                    16'hF192: data_out = 8'h83;
                    16'hF193: data_out = 8'h84;
                    16'hF194: data_out = 8'h85;
                    16'hF195: data_out = 8'h86;
                    16'hF196: data_out = 8'h87;
                    16'hF197: data_out = 8'h88;
                    16'hF198: data_out = 8'h89;
                    16'hF199: data_out = 8'h8A;
                    16'hF19A: data_out = 8'h8B;
                    16'hF19B: data_out = 8'h8C;
                    16'hF19C: data_out = 8'h8D;
                    16'hF19D: data_out = 8'h8E;
                    16'hF19E: data_out = 8'h8F;
                    16'hF19F: data_out = 8'h90;
                    16'hF1A0: data_out = 8'h91;
                    16'hF1A1: data_out = 8'h92;
                    16'hF1A2: data_out = 8'h93;
                    16'hF1A3: data_out = 8'h94;
                    16'hF1A4: data_out = 8'h95;
                    16'hF1A5: data_out = 8'h96;
                    16'hF1A6: data_out = 8'h97;
                    16'hF1A7: data_out = 8'h98;
                    16'hF1A8: data_out = 8'h99;
                    16'hF1A9: data_out = 8'h9A;
                    16'hF1AA: data_out = 8'h9B;
                    16'hF1AB: data_out = 8'h9C;
                    16'hF1AC: data_out = 8'h9D;
                    16'hF1AD: data_out = 8'h9E;
                    16'hF1AE: data_out = 8'h9F;
                    16'hF1AF: data_out = 8'hA0;
                    16'hF1B0: data_out = 8'hA1;
                    16'hF1B1: data_out = 8'hA2;
                    16'hF1B2: data_out = 8'hA3;
                    16'hF1B3: data_out = 8'hA4;
                    16'hF1B4: data_out = 8'hA5;
                    16'hF1B5: data_out = 8'hA6;
                    16'hF1B6: data_out = 8'hA7;
                    16'hF1B7: data_out = 8'hA8;
                    16'hF1B8: data_out = 8'hA9;
                    16'hF1B9: data_out = 8'hAA;
                    16'hF1BA: data_out = 8'hAB;
                    16'hF1BB: data_out = 8'hAC;
                    16'hF1BC: data_out = 8'hAD;
                    16'hF1BD: data_out = 8'hAE;
                    16'hF1BE: data_out = 8'hAF;
                    16'hF1BF: data_out = 8'hB0;
                    16'hF1C0: data_out = 8'hB1;
                    16'hF1C1: data_out = 8'hB2;
                    16'hF1C2: data_out = 8'hB3;
                    16'hF1C3: data_out = 8'hB4;
                    16'hF1C4: data_out = 8'hB5;
                    16'hF1C5: data_out = 8'hB6;
                    16'hF1C6: data_out = 8'hB7;
                    16'hF1C7: data_out = 8'hB8;
                    16'hF1C8: data_out = 8'hB9;
                    16'hF1C9: data_out = 8'hBA;
                    16'hF1CA: data_out = 8'hBB;
                    16'hF1CB: data_out = 8'hBC;
                    16'hF1CC: data_out = 8'hBD;
                    16'hF1CD: data_out = 8'hBE;
                    16'hF1CE: data_out = 8'hBF;
                    16'hF1CF: data_out = 8'hC0;
                    16'hF1D0: data_out = 8'hC1;
                    16'hF1D1: data_out = 8'hC2;
                    16'hF1D2: data_out = 8'hC3;
                    16'hF1D3: data_out = 8'hC4;
                    16'hF1D4: data_out = 8'hC5;
                    16'hF1D5: data_out = 8'hC6;
                    16'hF1D6: data_out = 8'hC7;
                    16'hF1D7: data_out = 8'hC8;
                    16'hF1D8: data_out = 8'hC9;
                    16'hF1D9: data_out = 8'hCA;
                    16'hF1DA: data_out = 8'hCB;
                    16'hF1DB: data_out = 8'hCC;
                    16'hF1DC: data_out = 8'hCD;
                    16'hF1DD: data_out = 8'hCE;
                    16'hF1DE: data_out = 8'hCF;
                    16'hF1DF: data_out = 8'hD0;
                    16'hF1E0: data_out = 8'hD1;
                    16'hF1E1: data_out = 8'hD2;
                    16'hF1E2: data_out = 8'hD3;
                    16'hF1E3: data_out = 8'hD4;
                    16'hF1E4: data_out = 8'hD5;
                    16'hF1E5: data_out = 8'hD6;
                    16'hF1E6: data_out = 8'hD7;
                    16'hF1E7: data_out = 8'hD8;
                    16'hF1E8: data_out = 8'hD9;
                    16'hF1E9: data_out = 8'hDA;
                    16'hF1EA: data_out = 8'hDB;
                    16'hF1EB: data_out = 8'hDC;
                    16'hF1EC: data_out = 8'hDD;
                    16'hF1ED: data_out = 8'hDE;
                    16'hF1EE: data_out = 8'hDF;
                    16'hF1EF: data_out = 8'hE0;
                    16'hF1F0: data_out = 8'hE1;
                    16'hF1F1: data_out = 8'hE2;
                    16'hF1F2: data_out = 8'hE3;
                    16'hF1F3: data_out = 8'hE4;
                    16'hF1F4: data_out = 8'hE5;
                    16'hF1F5: data_out = 8'hE6;
                    16'hF1F6: data_out = 8'hE7;
                    16'hF1F7: data_out = 8'hE8;
                    16'hF1F8: data_out = 8'hE9;
                    16'hF1F9: data_out = 8'hEA;
                    16'hF1FA: data_out = 8'hEB;
                    16'hF1FB: data_out = 8'hEC;
                    16'hF1FC: data_out = 8'hED;
                    16'hF1FD: data_out = 8'hEE;
                    16'hF1FE: data_out = 8'hEF;
                    16'hF1FF: data_out = 8'hF0;
                    16'hF200: data_out = 8'hF2;
                    16'hF201: data_out = 8'hF1;
                    16'hF202: data_out = 8'hF0;
                    16'hF203: data_out = 8'hEF;
                    16'hF204: data_out = 8'hEE;
                    16'hF205: data_out = 8'hED;
                    16'hF206: data_out = 8'hEC;
                    16'hF207: data_out = 8'hEB;
                    16'hF208: data_out = 8'hEA;
                    16'hF209: data_out = 8'hE9;
                    16'hF20A: data_out = 8'hE8;
                    16'hF20B: data_out = 8'hE7;
                    16'hF20C: data_out = 8'hE6;
                    16'hF20D: data_out = 8'hE5;
                    16'hF20E: data_out = 8'hE4;
                    16'hF20F: data_out = 8'hE3;
                    16'hF210: data_out = 8'hE2;
                    16'hF211: data_out = 8'hE1;
                    16'hF212: data_out = 8'hE0;
                    16'hF213: data_out = 8'hDF;
                    16'hF214: data_out = 8'hDE;
                    16'hF215: data_out = 8'hDD;
                    16'hF216: data_out = 8'hDC;
                    16'hF217: data_out = 8'hDB;
                    16'hF218: data_out = 8'hDA;
                    16'hF219: data_out = 8'hD9;
                    16'hF21A: data_out = 8'hD8;
                    16'hF21B: data_out = 8'hD7;
                    16'hF21C: data_out = 8'hD6;
                    16'hF21D: data_out = 8'hD5;
                    16'hF21E: data_out = 8'hD4;
                    16'hF21F: data_out = 8'hD3;
                    16'hF220: data_out = 8'hD2;
                    16'hF221: data_out = 8'hD1;
                    16'hF222: data_out = 8'hD0;
                    16'hF223: data_out = 8'hCF;
                    16'hF224: data_out = 8'hCE;
                    16'hF225: data_out = 8'hCD;
                    16'hF226: data_out = 8'hCC;
                    16'hF227: data_out = 8'hCB;
                    16'hF228: data_out = 8'hCA;
                    16'hF229: data_out = 8'hC9;
                    16'hF22A: data_out = 8'hC8;
                    16'hF22B: data_out = 8'hC7;
                    16'hF22C: data_out = 8'hC6;
                    16'hF22D: data_out = 8'hC5;
                    16'hF22E: data_out = 8'hC4;
                    16'hF22F: data_out = 8'hC3;
                    16'hF230: data_out = 8'hC2;
                    16'hF231: data_out = 8'hC1;
                    16'hF232: data_out = 8'hC0;
                    16'hF233: data_out = 8'hBF;
                    16'hF234: data_out = 8'hBE;
                    16'hF235: data_out = 8'hBD;
                    16'hF236: data_out = 8'hBC;
                    16'hF237: data_out = 8'hBB;
                    16'hF238: data_out = 8'hBA;
                    16'hF239: data_out = 8'hB9;
                    16'hF23A: data_out = 8'hB8;
                    16'hF23B: data_out = 8'hB7;
                    16'hF23C: data_out = 8'hB6;
                    16'hF23D: data_out = 8'hB5;
                    16'hF23E: data_out = 8'hB4;
                    16'hF23F: data_out = 8'hB3;
                    16'hF240: data_out = 8'hB2;
                    16'hF241: data_out = 8'hB1;
                    16'hF242: data_out = 8'hB0;
                    16'hF243: data_out = 8'hAF;
                    16'hF244: data_out = 8'hAE;
                    16'hF245: data_out = 8'hAD;
                    16'hF246: data_out = 8'hAC;
                    16'hF247: data_out = 8'hAB;
                    16'hF248: data_out = 8'hAA;
                    16'hF249: data_out = 8'hA9;
                    16'hF24A: data_out = 8'hA8;
                    16'hF24B: data_out = 8'hA7;
                    16'hF24C: data_out = 8'hA6;
                    16'hF24D: data_out = 8'hA5;
                    16'hF24E: data_out = 8'hA4;
                    16'hF24F: data_out = 8'hA3;
                    16'hF250: data_out = 8'hA2;
                    16'hF251: data_out = 8'hA1;
                    16'hF252: data_out = 8'hA0;
                    16'hF253: data_out = 8'h9F;
                    16'hF254: data_out = 8'h9E;
                    16'hF255: data_out = 8'h9D;
                    16'hF256: data_out = 8'h9C;
                    16'hF257: data_out = 8'h9B;
                    16'hF258: data_out = 8'h9A;
                    16'hF259: data_out = 8'h99;
                    16'hF25A: data_out = 8'h98;
                    16'hF25B: data_out = 8'h97;
                    16'hF25C: data_out = 8'h96;
                    16'hF25D: data_out = 8'h95;
                    16'hF25E: data_out = 8'h94;
                    16'hF25F: data_out = 8'h93;
                    16'hF260: data_out = 8'h92;
                    16'hF261: data_out = 8'h91;
                    16'hF262: data_out = 8'h90;
                    16'hF263: data_out = 8'h8F;
                    16'hF264: data_out = 8'h8E;
                    16'hF265: data_out = 8'h8D;
                    16'hF266: data_out = 8'h8C;
                    16'hF267: data_out = 8'h8B;
                    16'hF268: data_out = 8'h8A;
                    16'hF269: data_out = 8'h89;
                    16'hF26A: data_out = 8'h88;
                    16'hF26B: data_out = 8'h87;
                    16'hF26C: data_out = 8'h86;
                    16'hF26D: data_out = 8'h85;
                    16'hF26E: data_out = 8'h84;
                    16'hF26F: data_out = 8'h83;
                    16'hF270: data_out = 8'h82;
                    16'hF271: data_out = 8'h81;
                    16'hF272: data_out = 8'h0;
                    16'hF273: data_out = 8'h1;
                    16'hF274: data_out = 8'h2;
                    16'hF275: data_out = 8'h3;
                    16'hF276: data_out = 8'h4;
                    16'hF277: data_out = 8'h5;
                    16'hF278: data_out = 8'h6;
                    16'hF279: data_out = 8'h7;
                    16'hF27A: data_out = 8'h8;
                    16'hF27B: data_out = 8'h9;
                    16'hF27C: data_out = 8'hA;
                    16'hF27D: data_out = 8'hB;
                    16'hF27E: data_out = 8'hC;
                    16'hF27F: data_out = 8'hD;
                    16'hF280: data_out = 8'hF2;
                    16'hF281: data_out = 8'hF3;
                    16'hF282: data_out = 8'hF4;
                    16'hF283: data_out = 8'hF5;
                    16'hF284: data_out = 8'hF6;
                    16'hF285: data_out = 8'hF7;
                    16'hF286: data_out = 8'hF8;
                    16'hF287: data_out = 8'hF9;
                    16'hF288: data_out = 8'hFA;
                    16'hF289: data_out = 8'hFB;
                    16'hF28A: data_out = 8'hFC;
                    16'hF28B: data_out = 8'hFD;
                    16'hF28C: data_out = 8'hFE;
                    16'hF28D: data_out = 8'hFF;
                    16'hF28E: data_out = 8'h80;
                    16'hF28F: data_out = 8'h81;
                    16'hF290: data_out = 8'h82;
                    16'hF291: data_out = 8'h83;
                    16'hF292: data_out = 8'h84;
                    16'hF293: data_out = 8'h85;
                    16'hF294: data_out = 8'h86;
                    16'hF295: data_out = 8'h87;
                    16'hF296: data_out = 8'h88;
                    16'hF297: data_out = 8'h89;
                    16'hF298: data_out = 8'h8A;
                    16'hF299: data_out = 8'h8B;
                    16'hF29A: data_out = 8'h8C;
                    16'hF29B: data_out = 8'h8D;
                    16'hF29C: data_out = 8'h8E;
                    16'hF29D: data_out = 8'h8F;
                    16'hF29E: data_out = 8'h90;
                    16'hF29F: data_out = 8'h91;
                    16'hF2A0: data_out = 8'h92;
                    16'hF2A1: data_out = 8'h93;
                    16'hF2A2: data_out = 8'h94;
                    16'hF2A3: data_out = 8'h95;
                    16'hF2A4: data_out = 8'h96;
                    16'hF2A5: data_out = 8'h97;
                    16'hF2A6: data_out = 8'h98;
                    16'hF2A7: data_out = 8'h99;
                    16'hF2A8: data_out = 8'h9A;
                    16'hF2A9: data_out = 8'h9B;
                    16'hF2AA: data_out = 8'h9C;
                    16'hF2AB: data_out = 8'h9D;
                    16'hF2AC: data_out = 8'h9E;
                    16'hF2AD: data_out = 8'h9F;
                    16'hF2AE: data_out = 8'hA0;
                    16'hF2AF: data_out = 8'hA1;
                    16'hF2B0: data_out = 8'hA2;
                    16'hF2B1: data_out = 8'hA3;
                    16'hF2B2: data_out = 8'hA4;
                    16'hF2B3: data_out = 8'hA5;
                    16'hF2B4: data_out = 8'hA6;
                    16'hF2B5: data_out = 8'hA7;
                    16'hF2B6: data_out = 8'hA8;
                    16'hF2B7: data_out = 8'hA9;
                    16'hF2B8: data_out = 8'hAA;
                    16'hF2B9: data_out = 8'hAB;
                    16'hF2BA: data_out = 8'hAC;
                    16'hF2BB: data_out = 8'hAD;
                    16'hF2BC: data_out = 8'hAE;
                    16'hF2BD: data_out = 8'hAF;
                    16'hF2BE: data_out = 8'hB0;
                    16'hF2BF: data_out = 8'hB1;
                    16'hF2C0: data_out = 8'hB2;
                    16'hF2C1: data_out = 8'hB3;
                    16'hF2C2: data_out = 8'hB4;
                    16'hF2C3: data_out = 8'hB5;
                    16'hF2C4: data_out = 8'hB6;
                    16'hF2C5: data_out = 8'hB7;
                    16'hF2C6: data_out = 8'hB8;
                    16'hF2C7: data_out = 8'hB9;
                    16'hF2C8: data_out = 8'hBA;
                    16'hF2C9: data_out = 8'hBB;
                    16'hF2CA: data_out = 8'hBC;
                    16'hF2CB: data_out = 8'hBD;
                    16'hF2CC: data_out = 8'hBE;
                    16'hF2CD: data_out = 8'hBF;
                    16'hF2CE: data_out = 8'hC0;
                    16'hF2CF: data_out = 8'hC1;
                    16'hF2D0: data_out = 8'hC2;
                    16'hF2D1: data_out = 8'hC3;
                    16'hF2D2: data_out = 8'hC4;
                    16'hF2D3: data_out = 8'hC5;
                    16'hF2D4: data_out = 8'hC6;
                    16'hF2D5: data_out = 8'hC7;
                    16'hF2D6: data_out = 8'hC8;
                    16'hF2D7: data_out = 8'hC9;
                    16'hF2D8: data_out = 8'hCA;
                    16'hF2D9: data_out = 8'hCB;
                    16'hF2DA: data_out = 8'hCC;
                    16'hF2DB: data_out = 8'hCD;
                    16'hF2DC: data_out = 8'hCE;
                    16'hF2DD: data_out = 8'hCF;
                    16'hF2DE: data_out = 8'hD0;
                    16'hF2DF: data_out = 8'hD1;
                    16'hF2E0: data_out = 8'hD2;
                    16'hF2E1: data_out = 8'hD3;
                    16'hF2E2: data_out = 8'hD4;
                    16'hF2E3: data_out = 8'hD5;
                    16'hF2E4: data_out = 8'hD6;
                    16'hF2E5: data_out = 8'hD7;
                    16'hF2E6: data_out = 8'hD8;
                    16'hF2E7: data_out = 8'hD9;
                    16'hF2E8: data_out = 8'hDA;
                    16'hF2E9: data_out = 8'hDB;
                    16'hF2EA: data_out = 8'hDC;
                    16'hF2EB: data_out = 8'hDD;
                    16'hF2EC: data_out = 8'hDE;
                    16'hF2ED: data_out = 8'hDF;
                    16'hF2EE: data_out = 8'hE0;
                    16'hF2EF: data_out = 8'hE1;
                    16'hF2F0: data_out = 8'hE2;
                    16'hF2F1: data_out = 8'hE3;
                    16'hF2F2: data_out = 8'hE4;
                    16'hF2F3: data_out = 8'hE5;
                    16'hF2F4: data_out = 8'hE6;
                    16'hF2F5: data_out = 8'hE7;
                    16'hF2F6: data_out = 8'hE8;
                    16'hF2F7: data_out = 8'hE9;
                    16'hF2F8: data_out = 8'hEA;
                    16'hF2F9: data_out = 8'hEB;
                    16'hF2FA: data_out = 8'hEC;
                    16'hF2FB: data_out = 8'hED;
                    16'hF2FC: data_out = 8'hEE;
                    16'hF2FD: data_out = 8'hEF;
                    16'hF2FE: data_out = 8'hF0;
                    16'hF2FF: data_out = 8'hF1;
                    16'hF300: data_out = 8'hF3;
                    16'hF301: data_out = 8'hF2;
                    16'hF302: data_out = 8'hF1;
                    16'hF303: data_out = 8'hF0;
                    16'hF304: data_out = 8'hEF;
                    16'hF305: data_out = 8'hEE;
                    16'hF306: data_out = 8'hED;
                    16'hF307: data_out = 8'hEC;
                    16'hF308: data_out = 8'hEB;
                    16'hF309: data_out = 8'hEA;
                    16'hF30A: data_out = 8'hE9;
                    16'hF30B: data_out = 8'hE8;
                    16'hF30C: data_out = 8'hE7;
                    16'hF30D: data_out = 8'hE6;
                    16'hF30E: data_out = 8'hE5;
                    16'hF30F: data_out = 8'hE4;
                    16'hF310: data_out = 8'hE3;
                    16'hF311: data_out = 8'hE2;
                    16'hF312: data_out = 8'hE1;
                    16'hF313: data_out = 8'hE0;
                    16'hF314: data_out = 8'hDF;
                    16'hF315: data_out = 8'hDE;
                    16'hF316: data_out = 8'hDD;
                    16'hF317: data_out = 8'hDC;
                    16'hF318: data_out = 8'hDB;
                    16'hF319: data_out = 8'hDA;
                    16'hF31A: data_out = 8'hD9;
                    16'hF31B: data_out = 8'hD8;
                    16'hF31C: data_out = 8'hD7;
                    16'hF31D: data_out = 8'hD6;
                    16'hF31E: data_out = 8'hD5;
                    16'hF31F: data_out = 8'hD4;
                    16'hF320: data_out = 8'hD3;
                    16'hF321: data_out = 8'hD2;
                    16'hF322: data_out = 8'hD1;
                    16'hF323: data_out = 8'hD0;
                    16'hF324: data_out = 8'hCF;
                    16'hF325: data_out = 8'hCE;
                    16'hF326: data_out = 8'hCD;
                    16'hF327: data_out = 8'hCC;
                    16'hF328: data_out = 8'hCB;
                    16'hF329: data_out = 8'hCA;
                    16'hF32A: data_out = 8'hC9;
                    16'hF32B: data_out = 8'hC8;
                    16'hF32C: data_out = 8'hC7;
                    16'hF32D: data_out = 8'hC6;
                    16'hF32E: data_out = 8'hC5;
                    16'hF32F: data_out = 8'hC4;
                    16'hF330: data_out = 8'hC3;
                    16'hF331: data_out = 8'hC2;
                    16'hF332: data_out = 8'hC1;
                    16'hF333: data_out = 8'hC0;
                    16'hF334: data_out = 8'hBF;
                    16'hF335: data_out = 8'hBE;
                    16'hF336: data_out = 8'hBD;
                    16'hF337: data_out = 8'hBC;
                    16'hF338: data_out = 8'hBB;
                    16'hF339: data_out = 8'hBA;
                    16'hF33A: data_out = 8'hB9;
                    16'hF33B: data_out = 8'hB8;
                    16'hF33C: data_out = 8'hB7;
                    16'hF33D: data_out = 8'hB6;
                    16'hF33E: data_out = 8'hB5;
                    16'hF33F: data_out = 8'hB4;
                    16'hF340: data_out = 8'hB3;
                    16'hF341: data_out = 8'hB2;
                    16'hF342: data_out = 8'hB1;
                    16'hF343: data_out = 8'hB0;
                    16'hF344: data_out = 8'hAF;
                    16'hF345: data_out = 8'hAE;
                    16'hF346: data_out = 8'hAD;
                    16'hF347: data_out = 8'hAC;
                    16'hF348: data_out = 8'hAB;
                    16'hF349: data_out = 8'hAA;
                    16'hF34A: data_out = 8'hA9;
                    16'hF34B: data_out = 8'hA8;
                    16'hF34C: data_out = 8'hA7;
                    16'hF34D: data_out = 8'hA6;
                    16'hF34E: data_out = 8'hA5;
                    16'hF34F: data_out = 8'hA4;
                    16'hF350: data_out = 8'hA3;
                    16'hF351: data_out = 8'hA2;
                    16'hF352: data_out = 8'hA1;
                    16'hF353: data_out = 8'hA0;
                    16'hF354: data_out = 8'h9F;
                    16'hF355: data_out = 8'h9E;
                    16'hF356: data_out = 8'h9D;
                    16'hF357: data_out = 8'h9C;
                    16'hF358: data_out = 8'h9B;
                    16'hF359: data_out = 8'h9A;
                    16'hF35A: data_out = 8'h99;
                    16'hF35B: data_out = 8'h98;
                    16'hF35C: data_out = 8'h97;
                    16'hF35D: data_out = 8'h96;
                    16'hF35E: data_out = 8'h95;
                    16'hF35F: data_out = 8'h94;
                    16'hF360: data_out = 8'h93;
                    16'hF361: data_out = 8'h92;
                    16'hF362: data_out = 8'h91;
                    16'hF363: data_out = 8'h90;
                    16'hF364: data_out = 8'h8F;
                    16'hF365: data_out = 8'h8E;
                    16'hF366: data_out = 8'h8D;
                    16'hF367: data_out = 8'h8C;
                    16'hF368: data_out = 8'h8B;
                    16'hF369: data_out = 8'h8A;
                    16'hF36A: data_out = 8'h89;
                    16'hF36B: data_out = 8'h88;
                    16'hF36C: data_out = 8'h87;
                    16'hF36D: data_out = 8'h86;
                    16'hF36E: data_out = 8'h85;
                    16'hF36F: data_out = 8'h84;
                    16'hF370: data_out = 8'h83;
                    16'hF371: data_out = 8'h82;
                    16'hF372: data_out = 8'h81;
                    16'hF373: data_out = 8'h0;
                    16'hF374: data_out = 8'h1;
                    16'hF375: data_out = 8'h2;
                    16'hF376: data_out = 8'h3;
                    16'hF377: data_out = 8'h4;
                    16'hF378: data_out = 8'h5;
                    16'hF379: data_out = 8'h6;
                    16'hF37A: data_out = 8'h7;
                    16'hF37B: data_out = 8'h8;
                    16'hF37C: data_out = 8'h9;
                    16'hF37D: data_out = 8'hA;
                    16'hF37E: data_out = 8'hB;
                    16'hF37F: data_out = 8'hC;
                    16'hF380: data_out = 8'hF3;
                    16'hF381: data_out = 8'hF4;
                    16'hF382: data_out = 8'hF5;
                    16'hF383: data_out = 8'hF6;
                    16'hF384: data_out = 8'hF7;
                    16'hF385: data_out = 8'hF8;
                    16'hF386: data_out = 8'hF9;
                    16'hF387: data_out = 8'hFA;
                    16'hF388: data_out = 8'hFB;
                    16'hF389: data_out = 8'hFC;
                    16'hF38A: data_out = 8'hFD;
                    16'hF38B: data_out = 8'hFE;
                    16'hF38C: data_out = 8'hFF;
                    16'hF38D: data_out = 8'h80;
                    16'hF38E: data_out = 8'h81;
                    16'hF38F: data_out = 8'h82;
                    16'hF390: data_out = 8'h83;
                    16'hF391: data_out = 8'h84;
                    16'hF392: data_out = 8'h85;
                    16'hF393: data_out = 8'h86;
                    16'hF394: data_out = 8'h87;
                    16'hF395: data_out = 8'h88;
                    16'hF396: data_out = 8'h89;
                    16'hF397: data_out = 8'h8A;
                    16'hF398: data_out = 8'h8B;
                    16'hF399: data_out = 8'h8C;
                    16'hF39A: data_out = 8'h8D;
                    16'hF39B: data_out = 8'h8E;
                    16'hF39C: data_out = 8'h8F;
                    16'hF39D: data_out = 8'h90;
                    16'hF39E: data_out = 8'h91;
                    16'hF39F: data_out = 8'h92;
                    16'hF3A0: data_out = 8'h93;
                    16'hF3A1: data_out = 8'h94;
                    16'hF3A2: data_out = 8'h95;
                    16'hF3A3: data_out = 8'h96;
                    16'hF3A4: data_out = 8'h97;
                    16'hF3A5: data_out = 8'h98;
                    16'hF3A6: data_out = 8'h99;
                    16'hF3A7: data_out = 8'h9A;
                    16'hF3A8: data_out = 8'h9B;
                    16'hF3A9: data_out = 8'h9C;
                    16'hF3AA: data_out = 8'h9D;
                    16'hF3AB: data_out = 8'h9E;
                    16'hF3AC: data_out = 8'h9F;
                    16'hF3AD: data_out = 8'hA0;
                    16'hF3AE: data_out = 8'hA1;
                    16'hF3AF: data_out = 8'hA2;
                    16'hF3B0: data_out = 8'hA3;
                    16'hF3B1: data_out = 8'hA4;
                    16'hF3B2: data_out = 8'hA5;
                    16'hF3B3: data_out = 8'hA6;
                    16'hF3B4: data_out = 8'hA7;
                    16'hF3B5: data_out = 8'hA8;
                    16'hF3B6: data_out = 8'hA9;
                    16'hF3B7: data_out = 8'hAA;
                    16'hF3B8: data_out = 8'hAB;
                    16'hF3B9: data_out = 8'hAC;
                    16'hF3BA: data_out = 8'hAD;
                    16'hF3BB: data_out = 8'hAE;
                    16'hF3BC: data_out = 8'hAF;
                    16'hF3BD: data_out = 8'hB0;
                    16'hF3BE: data_out = 8'hB1;
                    16'hF3BF: data_out = 8'hB2;
                    16'hF3C0: data_out = 8'hB3;
                    16'hF3C1: data_out = 8'hB4;
                    16'hF3C2: data_out = 8'hB5;
                    16'hF3C3: data_out = 8'hB6;
                    16'hF3C4: data_out = 8'hB7;
                    16'hF3C5: data_out = 8'hB8;
                    16'hF3C6: data_out = 8'hB9;
                    16'hF3C7: data_out = 8'hBA;
                    16'hF3C8: data_out = 8'hBB;
                    16'hF3C9: data_out = 8'hBC;
                    16'hF3CA: data_out = 8'hBD;
                    16'hF3CB: data_out = 8'hBE;
                    16'hF3CC: data_out = 8'hBF;
                    16'hF3CD: data_out = 8'hC0;
                    16'hF3CE: data_out = 8'hC1;
                    16'hF3CF: data_out = 8'hC2;
                    16'hF3D0: data_out = 8'hC3;
                    16'hF3D1: data_out = 8'hC4;
                    16'hF3D2: data_out = 8'hC5;
                    16'hF3D3: data_out = 8'hC6;
                    16'hF3D4: data_out = 8'hC7;
                    16'hF3D5: data_out = 8'hC8;
                    16'hF3D6: data_out = 8'hC9;
                    16'hF3D7: data_out = 8'hCA;
                    16'hF3D8: data_out = 8'hCB;
                    16'hF3D9: data_out = 8'hCC;
                    16'hF3DA: data_out = 8'hCD;
                    16'hF3DB: data_out = 8'hCE;
                    16'hF3DC: data_out = 8'hCF;
                    16'hF3DD: data_out = 8'hD0;
                    16'hF3DE: data_out = 8'hD1;
                    16'hF3DF: data_out = 8'hD2;
                    16'hF3E0: data_out = 8'hD3;
                    16'hF3E1: data_out = 8'hD4;
                    16'hF3E2: data_out = 8'hD5;
                    16'hF3E3: data_out = 8'hD6;
                    16'hF3E4: data_out = 8'hD7;
                    16'hF3E5: data_out = 8'hD8;
                    16'hF3E6: data_out = 8'hD9;
                    16'hF3E7: data_out = 8'hDA;
                    16'hF3E8: data_out = 8'hDB;
                    16'hF3E9: data_out = 8'hDC;
                    16'hF3EA: data_out = 8'hDD;
                    16'hF3EB: data_out = 8'hDE;
                    16'hF3EC: data_out = 8'hDF;
                    16'hF3ED: data_out = 8'hE0;
                    16'hF3EE: data_out = 8'hE1;
                    16'hF3EF: data_out = 8'hE2;
                    16'hF3F0: data_out = 8'hE3;
                    16'hF3F1: data_out = 8'hE4;
                    16'hF3F2: data_out = 8'hE5;
                    16'hF3F3: data_out = 8'hE6;
                    16'hF3F4: data_out = 8'hE7;
                    16'hF3F5: data_out = 8'hE8;
                    16'hF3F6: data_out = 8'hE9;
                    16'hF3F7: data_out = 8'hEA;
                    16'hF3F8: data_out = 8'hEB;
                    16'hF3F9: data_out = 8'hEC;
                    16'hF3FA: data_out = 8'hED;
                    16'hF3FB: data_out = 8'hEE;
                    16'hF3FC: data_out = 8'hEF;
                    16'hF3FD: data_out = 8'hF0;
                    16'hF3FE: data_out = 8'hF1;
                    16'hF3FF: data_out = 8'hF2;
                    16'hF400: data_out = 8'hF4;
                    16'hF401: data_out = 8'hF3;
                    16'hF402: data_out = 8'hF2;
                    16'hF403: data_out = 8'hF1;
                    16'hF404: data_out = 8'hF0;
                    16'hF405: data_out = 8'hEF;
                    16'hF406: data_out = 8'hEE;
                    16'hF407: data_out = 8'hED;
                    16'hF408: data_out = 8'hEC;
                    16'hF409: data_out = 8'hEB;
                    16'hF40A: data_out = 8'hEA;
                    16'hF40B: data_out = 8'hE9;
                    16'hF40C: data_out = 8'hE8;
                    16'hF40D: data_out = 8'hE7;
                    16'hF40E: data_out = 8'hE6;
                    16'hF40F: data_out = 8'hE5;
                    16'hF410: data_out = 8'hE4;
                    16'hF411: data_out = 8'hE3;
                    16'hF412: data_out = 8'hE2;
                    16'hF413: data_out = 8'hE1;
                    16'hF414: data_out = 8'hE0;
                    16'hF415: data_out = 8'hDF;
                    16'hF416: data_out = 8'hDE;
                    16'hF417: data_out = 8'hDD;
                    16'hF418: data_out = 8'hDC;
                    16'hF419: data_out = 8'hDB;
                    16'hF41A: data_out = 8'hDA;
                    16'hF41B: data_out = 8'hD9;
                    16'hF41C: data_out = 8'hD8;
                    16'hF41D: data_out = 8'hD7;
                    16'hF41E: data_out = 8'hD6;
                    16'hF41F: data_out = 8'hD5;
                    16'hF420: data_out = 8'hD4;
                    16'hF421: data_out = 8'hD3;
                    16'hF422: data_out = 8'hD2;
                    16'hF423: data_out = 8'hD1;
                    16'hF424: data_out = 8'hD0;
                    16'hF425: data_out = 8'hCF;
                    16'hF426: data_out = 8'hCE;
                    16'hF427: data_out = 8'hCD;
                    16'hF428: data_out = 8'hCC;
                    16'hF429: data_out = 8'hCB;
                    16'hF42A: data_out = 8'hCA;
                    16'hF42B: data_out = 8'hC9;
                    16'hF42C: data_out = 8'hC8;
                    16'hF42D: data_out = 8'hC7;
                    16'hF42E: data_out = 8'hC6;
                    16'hF42F: data_out = 8'hC5;
                    16'hF430: data_out = 8'hC4;
                    16'hF431: data_out = 8'hC3;
                    16'hF432: data_out = 8'hC2;
                    16'hF433: data_out = 8'hC1;
                    16'hF434: data_out = 8'hC0;
                    16'hF435: data_out = 8'hBF;
                    16'hF436: data_out = 8'hBE;
                    16'hF437: data_out = 8'hBD;
                    16'hF438: data_out = 8'hBC;
                    16'hF439: data_out = 8'hBB;
                    16'hF43A: data_out = 8'hBA;
                    16'hF43B: data_out = 8'hB9;
                    16'hF43C: data_out = 8'hB8;
                    16'hF43D: data_out = 8'hB7;
                    16'hF43E: data_out = 8'hB6;
                    16'hF43F: data_out = 8'hB5;
                    16'hF440: data_out = 8'hB4;
                    16'hF441: data_out = 8'hB3;
                    16'hF442: data_out = 8'hB2;
                    16'hF443: data_out = 8'hB1;
                    16'hF444: data_out = 8'hB0;
                    16'hF445: data_out = 8'hAF;
                    16'hF446: data_out = 8'hAE;
                    16'hF447: data_out = 8'hAD;
                    16'hF448: data_out = 8'hAC;
                    16'hF449: data_out = 8'hAB;
                    16'hF44A: data_out = 8'hAA;
                    16'hF44B: data_out = 8'hA9;
                    16'hF44C: data_out = 8'hA8;
                    16'hF44D: data_out = 8'hA7;
                    16'hF44E: data_out = 8'hA6;
                    16'hF44F: data_out = 8'hA5;
                    16'hF450: data_out = 8'hA4;
                    16'hF451: data_out = 8'hA3;
                    16'hF452: data_out = 8'hA2;
                    16'hF453: data_out = 8'hA1;
                    16'hF454: data_out = 8'hA0;
                    16'hF455: data_out = 8'h9F;
                    16'hF456: data_out = 8'h9E;
                    16'hF457: data_out = 8'h9D;
                    16'hF458: data_out = 8'h9C;
                    16'hF459: data_out = 8'h9B;
                    16'hF45A: data_out = 8'h9A;
                    16'hF45B: data_out = 8'h99;
                    16'hF45C: data_out = 8'h98;
                    16'hF45D: data_out = 8'h97;
                    16'hF45E: data_out = 8'h96;
                    16'hF45F: data_out = 8'h95;
                    16'hF460: data_out = 8'h94;
                    16'hF461: data_out = 8'h93;
                    16'hF462: data_out = 8'h92;
                    16'hF463: data_out = 8'h91;
                    16'hF464: data_out = 8'h90;
                    16'hF465: data_out = 8'h8F;
                    16'hF466: data_out = 8'h8E;
                    16'hF467: data_out = 8'h8D;
                    16'hF468: data_out = 8'h8C;
                    16'hF469: data_out = 8'h8B;
                    16'hF46A: data_out = 8'h8A;
                    16'hF46B: data_out = 8'h89;
                    16'hF46C: data_out = 8'h88;
                    16'hF46D: data_out = 8'h87;
                    16'hF46E: data_out = 8'h86;
                    16'hF46F: data_out = 8'h85;
                    16'hF470: data_out = 8'h84;
                    16'hF471: data_out = 8'h83;
                    16'hF472: data_out = 8'h82;
                    16'hF473: data_out = 8'h81;
                    16'hF474: data_out = 8'h0;
                    16'hF475: data_out = 8'h1;
                    16'hF476: data_out = 8'h2;
                    16'hF477: data_out = 8'h3;
                    16'hF478: data_out = 8'h4;
                    16'hF479: data_out = 8'h5;
                    16'hF47A: data_out = 8'h6;
                    16'hF47B: data_out = 8'h7;
                    16'hF47C: data_out = 8'h8;
                    16'hF47D: data_out = 8'h9;
                    16'hF47E: data_out = 8'hA;
                    16'hF47F: data_out = 8'hB;
                    16'hF480: data_out = 8'hF4;
                    16'hF481: data_out = 8'hF5;
                    16'hF482: data_out = 8'hF6;
                    16'hF483: data_out = 8'hF7;
                    16'hF484: data_out = 8'hF8;
                    16'hF485: data_out = 8'hF9;
                    16'hF486: data_out = 8'hFA;
                    16'hF487: data_out = 8'hFB;
                    16'hF488: data_out = 8'hFC;
                    16'hF489: data_out = 8'hFD;
                    16'hF48A: data_out = 8'hFE;
                    16'hF48B: data_out = 8'hFF;
                    16'hF48C: data_out = 8'h80;
                    16'hF48D: data_out = 8'h81;
                    16'hF48E: data_out = 8'h82;
                    16'hF48F: data_out = 8'h83;
                    16'hF490: data_out = 8'h84;
                    16'hF491: data_out = 8'h85;
                    16'hF492: data_out = 8'h86;
                    16'hF493: data_out = 8'h87;
                    16'hF494: data_out = 8'h88;
                    16'hF495: data_out = 8'h89;
                    16'hF496: data_out = 8'h8A;
                    16'hF497: data_out = 8'h8B;
                    16'hF498: data_out = 8'h8C;
                    16'hF499: data_out = 8'h8D;
                    16'hF49A: data_out = 8'h8E;
                    16'hF49B: data_out = 8'h8F;
                    16'hF49C: data_out = 8'h90;
                    16'hF49D: data_out = 8'h91;
                    16'hF49E: data_out = 8'h92;
                    16'hF49F: data_out = 8'h93;
                    16'hF4A0: data_out = 8'h94;
                    16'hF4A1: data_out = 8'h95;
                    16'hF4A2: data_out = 8'h96;
                    16'hF4A3: data_out = 8'h97;
                    16'hF4A4: data_out = 8'h98;
                    16'hF4A5: data_out = 8'h99;
                    16'hF4A6: data_out = 8'h9A;
                    16'hF4A7: data_out = 8'h9B;
                    16'hF4A8: data_out = 8'h9C;
                    16'hF4A9: data_out = 8'h9D;
                    16'hF4AA: data_out = 8'h9E;
                    16'hF4AB: data_out = 8'h9F;
                    16'hF4AC: data_out = 8'hA0;
                    16'hF4AD: data_out = 8'hA1;
                    16'hF4AE: data_out = 8'hA2;
                    16'hF4AF: data_out = 8'hA3;
                    16'hF4B0: data_out = 8'hA4;
                    16'hF4B1: data_out = 8'hA5;
                    16'hF4B2: data_out = 8'hA6;
                    16'hF4B3: data_out = 8'hA7;
                    16'hF4B4: data_out = 8'hA8;
                    16'hF4B5: data_out = 8'hA9;
                    16'hF4B6: data_out = 8'hAA;
                    16'hF4B7: data_out = 8'hAB;
                    16'hF4B8: data_out = 8'hAC;
                    16'hF4B9: data_out = 8'hAD;
                    16'hF4BA: data_out = 8'hAE;
                    16'hF4BB: data_out = 8'hAF;
                    16'hF4BC: data_out = 8'hB0;
                    16'hF4BD: data_out = 8'hB1;
                    16'hF4BE: data_out = 8'hB2;
                    16'hF4BF: data_out = 8'hB3;
                    16'hF4C0: data_out = 8'hB4;
                    16'hF4C1: data_out = 8'hB5;
                    16'hF4C2: data_out = 8'hB6;
                    16'hF4C3: data_out = 8'hB7;
                    16'hF4C4: data_out = 8'hB8;
                    16'hF4C5: data_out = 8'hB9;
                    16'hF4C6: data_out = 8'hBA;
                    16'hF4C7: data_out = 8'hBB;
                    16'hF4C8: data_out = 8'hBC;
                    16'hF4C9: data_out = 8'hBD;
                    16'hF4CA: data_out = 8'hBE;
                    16'hF4CB: data_out = 8'hBF;
                    16'hF4CC: data_out = 8'hC0;
                    16'hF4CD: data_out = 8'hC1;
                    16'hF4CE: data_out = 8'hC2;
                    16'hF4CF: data_out = 8'hC3;
                    16'hF4D0: data_out = 8'hC4;
                    16'hF4D1: data_out = 8'hC5;
                    16'hF4D2: data_out = 8'hC6;
                    16'hF4D3: data_out = 8'hC7;
                    16'hF4D4: data_out = 8'hC8;
                    16'hF4D5: data_out = 8'hC9;
                    16'hF4D6: data_out = 8'hCA;
                    16'hF4D7: data_out = 8'hCB;
                    16'hF4D8: data_out = 8'hCC;
                    16'hF4D9: data_out = 8'hCD;
                    16'hF4DA: data_out = 8'hCE;
                    16'hF4DB: data_out = 8'hCF;
                    16'hF4DC: data_out = 8'hD0;
                    16'hF4DD: data_out = 8'hD1;
                    16'hF4DE: data_out = 8'hD2;
                    16'hF4DF: data_out = 8'hD3;
                    16'hF4E0: data_out = 8'hD4;
                    16'hF4E1: data_out = 8'hD5;
                    16'hF4E2: data_out = 8'hD6;
                    16'hF4E3: data_out = 8'hD7;
                    16'hF4E4: data_out = 8'hD8;
                    16'hF4E5: data_out = 8'hD9;
                    16'hF4E6: data_out = 8'hDA;
                    16'hF4E7: data_out = 8'hDB;
                    16'hF4E8: data_out = 8'hDC;
                    16'hF4E9: data_out = 8'hDD;
                    16'hF4EA: data_out = 8'hDE;
                    16'hF4EB: data_out = 8'hDF;
                    16'hF4EC: data_out = 8'hE0;
                    16'hF4ED: data_out = 8'hE1;
                    16'hF4EE: data_out = 8'hE2;
                    16'hF4EF: data_out = 8'hE3;
                    16'hF4F0: data_out = 8'hE4;
                    16'hF4F1: data_out = 8'hE5;
                    16'hF4F2: data_out = 8'hE6;
                    16'hF4F3: data_out = 8'hE7;
                    16'hF4F4: data_out = 8'hE8;
                    16'hF4F5: data_out = 8'hE9;
                    16'hF4F6: data_out = 8'hEA;
                    16'hF4F7: data_out = 8'hEB;
                    16'hF4F8: data_out = 8'hEC;
                    16'hF4F9: data_out = 8'hED;
                    16'hF4FA: data_out = 8'hEE;
                    16'hF4FB: data_out = 8'hEF;
                    16'hF4FC: data_out = 8'hF0;
                    16'hF4FD: data_out = 8'hF1;
                    16'hF4FE: data_out = 8'hF2;
                    16'hF4FF: data_out = 8'hF3;
                    16'hF500: data_out = 8'hF5;
                    16'hF501: data_out = 8'hF4;
                    16'hF502: data_out = 8'hF3;
                    16'hF503: data_out = 8'hF2;
                    16'hF504: data_out = 8'hF1;
                    16'hF505: data_out = 8'hF0;
                    16'hF506: data_out = 8'hEF;
                    16'hF507: data_out = 8'hEE;
                    16'hF508: data_out = 8'hED;
                    16'hF509: data_out = 8'hEC;
                    16'hF50A: data_out = 8'hEB;
                    16'hF50B: data_out = 8'hEA;
                    16'hF50C: data_out = 8'hE9;
                    16'hF50D: data_out = 8'hE8;
                    16'hF50E: data_out = 8'hE7;
                    16'hF50F: data_out = 8'hE6;
                    16'hF510: data_out = 8'hE5;
                    16'hF511: data_out = 8'hE4;
                    16'hF512: data_out = 8'hE3;
                    16'hF513: data_out = 8'hE2;
                    16'hF514: data_out = 8'hE1;
                    16'hF515: data_out = 8'hE0;
                    16'hF516: data_out = 8'hDF;
                    16'hF517: data_out = 8'hDE;
                    16'hF518: data_out = 8'hDD;
                    16'hF519: data_out = 8'hDC;
                    16'hF51A: data_out = 8'hDB;
                    16'hF51B: data_out = 8'hDA;
                    16'hF51C: data_out = 8'hD9;
                    16'hF51D: data_out = 8'hD8;
                    16'hF51E: data_out = 8'hD7;
                    16'hF51F: data_out = 8'hD6;
                    16'hF520: data_out = 8'hD5;
                    16'hF521: data_out = 8'hD4;
                    16'hF522: data_out = 8'hD3;
                    16'hF523: data_out = 8'hD2;
                    16'hF524: data_out = 8'hD1;
                    16'hF525: data_out = 8'hD0;
                    16'hF526: data_out = 8'hCF;
                    16'hF527: data_out = 8'hCE;
                    16'hF528: data_out = 8'hCD;
                    16'hF529: data_out = 8'hCC;
                    16'hF52A: data_out = 8'hCB;
                    16'hF52B: data_out = 8'hCA;
                    16'hF52C: data_out = 8'hC9;
                    16'hF52D: data_out = 8'hC8;
                    16'hF52E: data_out = 8'hC7;
                    16'hF52F: data_out = 8'hC6;
                    16'hF530: data_out = 8'hC5;
                    16'hF531: data_out = 8'hC4;
                    16'hF532: data_out = 8'hC3;
                    16'hF533: data_out = 8'hC2;
                    16'hF534: data_out = 8'hC1;
                    16'hF535: data_out = 8'hC0;
                    16'hF536: data_out = 8'hBF;
                    16'hF537: data_out = 8'hBE;
                    16'hF538: data_out = 8'hBD;
                    16'hF539: data_out = 8'hBC;
                    16'hF53A: data_out = 8'hBB;
                    16'hF53B: data_out = 8'hBA;
                    16'hF53C: data_out = 8'hB9;
                    16'hF53D: data_out = 8'hB8;
                    16'hF53E: data_out = 8'hB7;
                    16'hF53F: data_out = 8'hB6;
                    16'hF540: data_out = 8'hB5;
                    16'hF541: data_out = 8'hB4;
                    16'hF542: data_out = 8'hB3;
                    16'hF543: data_out = 8'hB2;
                    16'hF544: data_out = 8'hB1;
                    16'hF545: data_out = 8'hB0;
                    16'hF546: data_out = 8'hAF;
                    16'hF547: data_out = 8'hAE;
                    16'hF548: data_out = 8'hAD;
                    16'hF549: data_out = 8'hAC;
                    16'hF54A: data_out = 8'hAB;
                    16'hF54B: data_out = 8'hAA;
                    16'hF54C: data_out = 8'hA9;
                    16'hF54D: data_out = 8'hA8;
                    16'hF54E: data_out = 8'hA7;
                    16'hF54F: data_out = 8'hA6;
                    16'hF550: data_out = 8'hA5;
                    16'hF551: data_out = 8'hA4;
                    16'hF552: data_out = 8'hA3;
                    16'hF553: data_out = 8'hA2;
                    16'hF554: data_out = 8'hA1;
                    16'hF555: data_out = 8'hA0;
                    16'hF556: data_out = 8'h9F;
                    16'hF557: data_out = 8'h9E;
                    16'hF558: data_out = 8'h9D;
                    16'hF559: data_out = 8'h9C;
                    16'hF55A: data_out = 8'h9B;
                    16'hF55B: data_out = 8'h9A;
                    16'hF55C: data_out = 8'h99;
                    16'hF55D: data_out = 8'h98;
                    16'hF55E: data_out = 8'h97;
                    16'hF55F: data_out = 8'h96;
                    16'hF560: data_out = 8'h95;
                    16'hF561: data_out = 8'h94;
                    16'hF562: data_out = 8'h93;
                    16'hF563: data_out = 8'h92;
                    16'hF564: data_out = 8'h91;
                    16'hF565: data_out = 8'h90;
                    16'hF566: data_out = 8'h8F;
                    16'hF567: data_out = 8'h8E;
                    16'hF568: data_out = 8'h8D;
                    16'hF569: data_out = 8'h8C;
                    16'hF56A: data_out = 8'h8B;
                    16'hF56B: data_out = 8'h8A;
                    16'hF56C: data_out = 8'h89;
                    16'hF56D: data_out = 8'h88;
                    16'hF56E: data_out = 8'h87;
                    16'hF56F: data_out = 8'h86;
                    16'hF570: data_out = 8'h85;
                    16'hF571: data_out = 8'h84;
                    16'hF572: data_out = 8'h83;
                    16'hF573: data_out = 8'h82;
                    16'hF574: data_out = 8'h81;
                    16'hF575: data_out = 8'h0;
                    16'hF576: data_out = 8'h1;
                    16'hF577: data_out = 8'h2;
                    16'hF578: data_out = 8'h3;
                    16'hF579: data_out = 8'h4;
                    16'hF57A: data_out = 8'h5;
                    16'hF57B: data_out = 8'h6;
                    16'hF57C: data_out = 8'h7;
                    16'hF57D: data_out = 8'h8;
                    16'hF57E: data_out = 8'h9;
                    16'hF57F: data_out = 8'hA;
                    16'hF580: data_out = 8'hF5;
                    16'hF581: data_out = 8'hF6;
                    16'hF582: data_out = 8'hF7;
                    16'hF583: data_out = 8'hF8;
                    16'hF584: data_out = 8'hF9;
                    16'hF585: data_out = 8'hFA;
                    16'hF586: data_out = 8'hFB;
                    16'hF587: data_out = 8'hFC;
                    16'hF588: data_out = 8'hFD;
                    16'hF589: data_out = 8'hFE;
                    16'hF58A: data_out = 8'hFF;
                    16'hF58B: data_out = 8'h80;
                    16'hF58C: data_out = 8'h81;
                    16'hF58D: data_out = 8'h82;
                    16'hF58E: data_out = 8'h83;
                    16'hF58F: data_out = 8'h84;
                    16'hF590: data_out = 8'h85;
                    16'hF591: data_out = 8'h86;
                    16'hF592: data_out = 8'h87;
                    16'hF593: data_out = 8'h88;
                    16'hF594: data_out = 8'h89;
                    16'hF595: data_out = 8'h8A;
                    16'hF596: data_out = 8'h8B;
                    16'hF597: data_out = 8'h8C;
                    16'hF598: data_out = 8'h8D;
                    16'hF599: data_out = 8'h8E;
                    16'hF59A: data_out = 8'h8F;
                    16'hF59B: data_out = 8'h90;
                    16'hF59C: data_out = 8'h91;
                    16'hF59D: data_out = 8'h92;
                    16'hF59E: data_out = 8'h93;
                    16'hF59F: data_out = 8'h94;
                    16'hF5A0: data_out = 8'h95;
                    16'hF5A1: data_out = 8'h96;
                    16'hF5A2: data_out = 8'h97;
                    16'hF5A3: data_out = 8'h98;
                    16'hF5A4: data_out = 8'h99;
                    16'hF5A5: data_out = 8'h9A;
                    16'hF5A6: data_out = 8'h9B;
                    16'hF5A7: data_out = 8'h9C;
                    16'hF5A8: data_out = 8'h9D;
                    16'hF5A9: data_out = 8'h9E;
                    16'hF5AA: data_out = 8'h9F;
                    16'hF5AB: data_out = 8'hA0;
                    16'hF5AC: data_out = 8'hA1;
                    16'hF5AD: data_out = 8'hA2;
                    16'hF5AE: data_out = 8'hA3;
                    16'hF5AF: data_out = 8'hA4;
                    16'hF5B0: data_out = 8'hA5;
                    16'hF5B1: data_out = 8'hA6;
                    16'hF5B2: data_out = 8'hA7;
                    16'hF5B3: data_out = 8'hA8;
                    16'hF5B4: data_out = 8'hA9;
                    16'hF5B5: data_out = 8'hAA;
                    16'hF5B6: data_out = 8'hAB;
                    16'hF5B7: data_out = 8'hAC;
                    16'hF5B8: data_out = 8'hAD;
                    16'hF5B9: data_out = 8'hAE;
                    16'hF5BA: data_out = 8'hAF;
                    16'hF5BB: data_out = 8'hB0;
                    16'hF5BC: data_out = 8'hB1;
                    16'hF5BD: data_out = 8'hB2;
                    16'hF5BE: data_out = 8'hB3;
                    16'hF5BF: data_out = 8'hB4;
                    16'hF5C0: data_out = 8'hB5;
                    16'hF5C1: data_out = 8'hB6;
                    16'hF5C2: data_out = 8'hB7;
                    16'hF5C3: data_out = 8'hB8;
                    16'hF5C4: data_out = 8'hB9;
                    16'hF5C5: data_out = 8'hBA;
                    16'hF5C6: data_out = 8'hBB;
                    16'hF5C7: data_out = 8'hBC;
                    16'hF5C8: data_out = 8'hBD;
                    16'hF5C9: data_out = 8'hBE;
                    16'hF5CA: data_out = 8'hBF;
                    16'hF5CB: data_out = 8'hC0;
                    16'hF5CC: data_out = 8'hC1;
                    16'hF5CD: data_out = 8'hC2;
                    16'hF5CE: data_out = 8'hC3;
                    16'hF5CF: data_out = 8'hC4;
                    16'hF5D0: data_out = 8'hC5;
                    16'hF5D1: data_out = 8'hC6;
                    16'hF5D2: data_out = 8'hC7;
                    16'hF5D3: data_out = 8'hC8;
                    16'hF5D4: data_out = 8'hC9;
                    16'hF5D5: data_out = 8'hCA;
                    16'hF5D6: data_out = 8'hCB;
                    16'hF5D7: data_out = 8'hCC;
                    16'hF5D8: data_out = 8'hCD;
                    16'hF5D9: data_out = 8'hCE;
                    16'hF5DA: data_out = 8'hCF;
                    16'hF5DB: data_out = 8'hD0;
                    16'hF5DC: data_out = 8'hD1;
                    16'hF5DD: data_out = 8'hD2;
                    16'hF5DE: data_out = 8'hD3;
                    16'hF5DF: data_out = 8'hD4;
                    16'hF5E0: data_out = 8'hD5;
                    16'hF5E1: data_out = 8'hD6;
                    16'hF5E2: data_out = 8'hD7;
                    16'hF5E3: data_out = 8'hD8;
                    16'hF5E4: data_out = 8'hD9;
                    16'hF5E5: data_out = 8'hDA;
                    16'hF5E6: data_out = 8'hDB;
                    16'hF5E7: data_out = 8'hDC;
                    16'hF5E8: data_out = 8'hDD;
                    16'hF5E9: data_out = 8'hDE;
                    16'hF5EA: data_out = 8'hDF;
                    16'hF5EB: data_out = 8'hE0;
                    16'hF5EC: data_out = 8'hE1;
                    16'hF5ED: data_out = 8'hE2;
                    16'hF5EE: data_out = 8'hE3;
                    16'hF5EF: data_out = 8'hE4;
                    16'hF5F0: data_out = 8'hE5;
                    16'hF5F1: data_out = 8'hE6;
                    16'hF5F2: data_out = 8'hE7;
                    16'hF5F3: data_out = 8'hE8;
                    16'hF5F4: data_out = 8'hE9;
                    16'hF5F5: data_out = 8'hEA;
                    16'hF5F6: data_out = 8'hEB;
                    16'hF5F7: data_out = 8'hEC;
                    16'hF5F8: data_out = 8'hED;
                    16'hF5F9: data_out = 8'hEE;
                    16'hF5FA: data_out = 8'hEF;
                    16'hF5FB: data_out = 8'hF0;
                    16'hF5FC: data_out = 8'hF1;
                    16'hF5FD: data_out = 8'hF2;
                    16'hF5FE: data_out = 8'hF3;
                    16'hF5FF: data_out = 8'hF4;
                    16'hF600: data_out = 8'hF6;
                    16'hF601: data_out = 8'hF5;
                    16'hF602: data_out = 8'hF4;
                    16'hF603: data_out = 8'hF3;
                    16'hF604: data_out = 8'hF2;
                    16'hF605: data_out = 8'hF1;
                    16'hF606: data_out = 8'hF0;
                    16'hF607: data_out = 8'hEF;
                    16'hF608: data_out = 8'hEE;
                    16'hF609: data_out = 8'hED;
                    16'hF60A: data_out = 8'hEC;
                    16'hF60B: data_out = 8'hEB;
                    16'hF60C: data_out = 8'hEA;
                    16'hF60D: data_out = 8'hE9;
                    16'hF60E: data_out = 8'hE8;
                    16'hF60F: data_out = 8'hE7;
                    16'hF610: data_out = 8'hE6;
                    16'hF611: data_out = 8'hE5;
                    16'hF612: data_out = 8'hE4;
                    16'hF613: data_out = 8'hE3;
                    16'hF614: data_out = 8'hE2;
                    16'hF615: data_out = 8'hE1;
                    16'hF616: data_out = 8'hE0;
                    16'hF617: data_out = 8'hDF;
                    16'hF618: data_out = 8'hDE;
                    16'hF619: data_out = 8'hDD;
                    16'hF61A: data_out = 8'hDC;
                    16'hF61B: data_out = 8'hDB;
                    16'hF61C: data_out = 8'hDA;
                    16'hF61D: data_out = 8'hD9;
                    16'hF61E: data_out = 8'hD8;
                    16'hF61F: data_out = 8'hD7;
                    16'hF620: data_out = 8'hD6;
                    16'hF621: data_out = 8'hD5;
                    16'hF622: data_out = 8'hD4;
                    16'hF623: data_out = 8'hD3;
                    16'hF624: data_out = 8'hD2;
                    16'hF625: data_out = 8'hD1;
                    16'hF626: data_out = 8'hD0;
                    16'hF627: data_out = 8'hCF;
                    16'hF628: data_out = 8'hCE;
                    16'hF629: data_out = 8'hCD;
                    16'hF62A: data_out = 8'hCC;
                    16'hF62B: data_out = 8'hCB;
                    16'hF62C: data_out = 8'hCA;
                    16'hF62D: data_out = 8'hC9;
                    16'hF62E: data_out = 8'hC8;
                    16'hF62F: data_out = 8'hC7;
                    16'hF630: data_out = 8'hC6;
                    16'hF631: data_out = 8'hC5;
                    16'hF632: data_out = 8'hC4;
                    16'hF633: data_out = 8'hC3;
                    16'hF634: data_out = 8'hC2;
                    16'hF635: data_out = 8'hC1;
                    16'hF636: data_out = 8'hC0;
                    16'hF637: data_out = 8'hBF;
                    16'hF638: data_out = 8'hBE;
                    16'hF639: data_out = 8'hBD;
                    16'hF63A: data_out = 8'hBC;
                    16'hF63B: data_out = 8'hBB;
                    16'hF63C: data_out = 8'hBA;
                    16'hF63D: data_out = 8'hB9;
                    16'hF63E: data_out = 8'hB8;
                    16'hF63F: data_out = 8'hB7;
                    16'hF640: data_out = 8'hB6;
                    16'hF641: data_out = 8'hB5;
                    16'hF642: data_out = 8'hB4;
                    16'hF643: data_out = 8'hB3;
                    16'hF644: data_out = 8'hB2;
                    16'hF645: data_out = 8'hB1;
                    16'hF646: data_out = 8'hB0;
                    16'hF647: data_out = 8'hAF;
                    16'hF648: data_out = 8'hAE;
                    16'hF649: data_out = 8'hAD;
                    16'hF64A: data_out = 8'hAC;
                    16'hF64B: data_out = 8'hAB;
                    16'hF64C: data_out = 8'hAA;
                    16'hF64D: data_out = 8'hA9;
                    16'hF64E: data_out = 8'hA8;
                    16'hF64F: data_out = 8'hA7;
                    16'hF650: data_out = 8'hA6;
                    16'hF651: data_out = 8'hA5;
                    16'hF652: data_out = 8'hA4;
                    16'hF653: data_out = 8'hA3;
                    16'hF654: data_out = 8'hA2;
                    16'hF655: data_out = 8'hA1;
                    16'hF656: data_out = 8'hA0;
                    16'hF657: data_out = 8'h9F;
                    16'hF658: data_out = 8'h9E;
                    16'hF659: data_out = 8'h9D;
                    16'hF65A: data_out = 8'h9C;
                    16'hF65B: data_out = 8'h9B;
                    16'hF65C: data_out = 8'h9A;
                    16'hF65D: data_out = 8'h99;
                    16'hF65E: data_out = 8'h98;
                    16'hF65F: data_out = 8'h97;
                    16'hF660: data_out = 8'h96;
                    16'hF661: data_out = 8'h95;
                    16'hF662: data_out = 8'h94;
                    16'hF663: data_out = 8'h93;
                    16'hF664: data_out = 8'h92;
                    16'hF665: data_out = 8'h91;
                    16'hF666: data_out = 8'h90;
                    16'hF667: data_out = 8'h8F;
                    16'hF668: data_out = 8'h8E;
                    16'hF669: data_out = 8'h8D;
                    16'hF66A: data_out = 8'h8C;
                    16'hF66B: data_out = 8'h8B;
                    16'hF66C: data_out = 8'h8A;
                    16'hF66D: data_out = 8'h89;
                    16'hF66E: data_out = 8'h88;
                    16'hF66F: data_out = 8'h87;
                    16'hF670: data_out = 8'h86;
                    16'hF671: data_out = 8'h85;
                    16'hF672: data_out = 8'h84;
                    16'hF673: data_out = 8'h83;
                    16'hF674: data_out = 8'h82;
                    16'hF675: data_out = 8'h81;
                    16'hF676: data_out = 8'h0;
                    16'hF677: data_out = 8'h1;
                    16'hF678: data_out = 8'h2;
                    16'hF679: data_out = 8'h3;
                    16'hF67A: data_out = 8'h4;
                    16'hF67B: data_out = 8'h5;
                    16'hF67C: data_out = 8'h6;
                    16'hF67D: data_out = 8'h7;
                    16'hF67E: data_out = 8'h8;
                    16'hF67F: data_out = 8'h9;
                    16'hF680: data_out = 8'hF6;
                    16'hF681: data_out = 8'hF7;
                    16'hF682: data_out = 8'hF8;
                    16'hF683: data_out = 8'hF9;
                    16'hF684: data_out = 8'hFA;
                    16'hF685: data_out = 8'hFB;
                    16'hF686: data_out = 8'hFC;
                    16'hF687: data_out = 8'hFD;
                    16'hF688: data_out = 8'hFE;
                    16'hF689: data_out = 8'hFF;
                    16'hF68A: data_out = 8'h80;
                    16'hF68B: data_out = 8'h81;
                    16'hF68C: data_out = 8'h82;
                    16'hF68D: data_out = 8'h83;
                    16'hF68E: data_out = 8'h84;
                    16'hF68F: data_out = 8'h85;
                    16'hF690: data_out = 8'h86;
                    16'hF691: data_out = 8'h87;
                    16'hF692: data_out = 8'h88;
                    16'hF693: data_out = 8'h89;
                    16'hF694: data_out = 8'h8A;
                    16'hF695: data_out = 8'h8B;
                    16'hF696: data_out = 8'h8C;
                    16'hF697: data_out = 8'h8D;
                    16'hF698: data_out = 8'h8E;
                    16'hF699: data_out = 8'h8F;
                    16'hF69A: data_out = 8'h90;
                    16'hF69B: data_out = 8'h91;
                    16'hF69C: data_out = 8'h92;
                    16'hF69D: data_out = 8'h93;
                    16'hF69E: data_out = 8'h94;
                    16'hF69F: data_out = 8'h95;
                    16'hF6A0: data_out = 8'h96;
                    16'hF6A1: data_out = 8'h97;
                    16'hF6A2: data_out = 8'h98;
                    16'hF6A3: data_out = 8'h99;
                    16'hF6A4: data_out = 8'h9A;
                    16'hF6A5: data_out = 8'h9B;
                    16'hF6A6: data_out = 8'h9C;
                    16'hF6A7: data_out = 8'h9D;
                    16'hF6A8: data_out = 8'h9E;
                    16'hF6A9: data_out = 8'h9F;
                    16'hF6AA: data_out = 8'hA0;
                    16'hF6AB: data_out = 8'hA1;
                    16'hF6AC: data_out = 8'hA2;
                    16'hF6AD: data_out = 8'hA3;
                    16'hF6AE: data_out = 8'hA4;
                    16'hF6AF: data_out = 8'hA5;
                    16'hF6B0: data_out = 8'hA6;
                    16'hF6B1: data_out = 8'hA7;
                    16'hF6B2: data_out = 8'hA8;
                    16'hF6B3: data_out = 8'hA9;
                    16'hF6B4: data_out = 8'hAA;
                    16'hF6B5: data_out = 8'hAB;
                    16'hF6B6: data_out = 8'hAC;
                    16'hF6B7: data_out = 8'hAD;
                    16'hF6B8: data_out = 8'hAE;
                    16'hF6B9: data_out = 8'hAF;
                    16'hF6BA: data_out = 8'hB0;
                    16'hF6BB: data_out = 8'hB1;
                    16'hF6BC: data_out = 8'hB2;
                    16'hF6BD: data_out = 8'hB3;
                    16'hF6BE: data_out = 8'hB4;
                    16'hF6BF: data_out = 8'hB5;
                    16'hF6C0: data_out = 8'hB6;
                    16'hF6C1: data_out = 8'hB7;
                    16'hF6C2: data_out = 8'hB8;
                    16'hF6C3: data_out = 8'hB9;
                    16'hF6C4: data_out = 8'hBA;
                    16'hF6C5: data_out = 8'hBB;
                    16'hF6C6: data_out = 8'hBC;
                    16'hF6C7: data_out = 8'hBD;
                    16'hF6C8: data_out = 8'hBE;
                    16'hF6C9: data_out = 8'hBF;
                    16'hF6CA: data_out = 8'hC0;
                    16'hF6CB: data_out = 8'hC1;
                    16'hF6CC: data_out = 8'hC2;
                    16'hF6CD: data_out = 8'hC3;
                    16'hF6CE: data_out = 8'hC4;
                    16'hF6CF: data_out = 8'hC5;
                    16'hF6D0: data_out = 8'hC6;
                    16'hF6D1: data_out = 8'hC7;
                    16'hF6D2: data_out = 8'hC8;
                    16'hF6D3: data_out = 8'hC9;
                    16'hF6D4: data_out = 8'hCA;
                    16'hF6D5: data_out = 8'hCB;
                    16'hF6D6: data_out = 8'hCC;
                    16'hF6D7: data_out = 8'hCD;
                    16'hF6D8: data_out = 8'hCE;
                    16'hF6D9: data_out = 8'hCF;
                    16'hF6DA: data_out = 8'hD0;
                    16'hF6DB: data_out = 8'hD1;
                    16'hF6DC: data_out = 8'hD2;
                    16'hF6DD: data_out = 8'hD3;
                    16'hF6DE: data_out = 8'hD4;
                    16'hF6DF: data_out = 8'hD5;
                    16'hF6E0: data_out = 8'hD6;
                    16'hF6E1: data_out = 8'hD7;
                    16'hF6E2: data_out = 8'hD8;
                    16'hF6E3: data_out = 8'hD9;
                    16'hF6E4: data_out = 8'hDA;
                    16'hF6E5: data_out = 8'hDB;
                    16'hF6E6: data_out = 8'hDC;
                    16'hF6E7: data_out = 8'hDD;
                    16'hF6E8: data_out = 8'hDE;
                    16'hF6E9: data_out = 8'hDF;
                    16'hF6EA: data_out = 8'hE0;
                    16'hF6EB: data_out = 8'hE1;
                    16'hF6EC: data_out = 8'hE2;
                    16'hF6ED: data_out = 8'hE3;
                    16'hF6EE: data_out = 8'hE4;
                    16'hF6EF: data_out = 8'hE5;
                    16'hF6F0: data_out = 8'hE6;
                    16'hF6F1: data_out = 8'hE7;
                    16'hF6F2: data_out = 8'hE8;
                    16'hF6F3: data_out = 8'hE9;
                    16'hF6F4: data_out = 8'hEA;
                    16'hF6F5: data_out = 8'hEB;
                    16'hF6F6: data_out = 8'hEC;
                    16'hF6F7: data_out = 8'hED;
                    16'hF6F8: data_out = 8'hEE;
                    16'hF6F9: data_out = 8'hEF;
                    16'hF6FA: data_out = 8'hF0;
                    16'hF6FB: data_out = 8'hF1;
                    16'hF6FC: data_out = 8'hF2;
                    16'hF6FD: data_out = 8'hF3;
                    16'hF6FE: data_out = 8'hF4;
                    16'hF6FF: data_out = 8'hF5;
                    16'hF700: data_out = 8'hF7;
                    16'hF701: data_out = 8'hF6;
                    16'hF702: data_out = 8'hF5;
                    16'hF703: data_out = 8'hF4;
                    16'hF704: data_out = 8'hF3;
                    16'hF705: data_out = 8'hF2;
                    16'hF706: data_out = 8'hF1;
                    16'hF707: data_out = 8'hF0;
                    16'hF708: data_out = 8'hEF;
                    16'hF709: data_out = 8'hEE;
                    16'hF70A: data_out = 8'hED;
                    16'hF70B: data_out = 8'hEC;
                    16'hF70C: data_out = 8'hEB;
                    16'hF70D: data_out = 8'hEA;
                    16'hF70E: data_out = 8'hE9;
                    16'hF70F: data_out = 8'hE8;
                    16'hF710: data_out = 8'hE7;
                    16'hF711: data_out = 8'hE6;
                    16'hF712: data_out = 8'hE5;
                    16'hF713: data_out = 8'hE4;
                    16'hF714: data_out = 8'hE3;
                    16'hF715: data_out = 8'hE2;
                    16'hF716: data_out = 8'hE1;
                    16'hF717: data_out = 8'hE0;
                    16'hF718: data_out = 8'hDF;
                    16'hF719: data_out = 8'hDE;
                    16'hF71A: data_out = 8'hDD;
                    16'hF71B: data_out = 8'hDC;
                    16'hF71C: data_out = 8'hDB;
                    16'hF71D: data_out = 8'hDA;
                    16'hF71E: data_out = 8'hD9;
                    16'hF71F: data_out = 8'hD8;
                    16'hF720: data_out = 8'hD7;
                    16'hF721: data_out = 8'hD6;
                    16'hF722: data_out = 8'hD5;
                    16'hF723: data_out = 8'hD4;
                    16'hF724: data_out = 8'hD3;
                    16'hF725: data_out = 8'hD2;
                    16'hF726: data_out = 8'hD1;
                    16'hF727: data_out = 8'hD0;
                    16'hF728: data_out = 8'hCF;
                    16'hF729: data_out = 8'hCE;
                    16'hF72A: data_out = 8'hCD;
                    16'hF72B: data_out = 8'hCC;
                    16'hF72C: data_out = 8'hCB;
                    16'hF72D: data_out = 8'hCA;
                    16'hF72E: data_out = 8'hC9;
                    16'hF72F: data_out = 8'hC8;
                    16'hF730: data_out = 8'hC7;
                    16'hF731: data_out = 8'hC6;
                    16'hF732: data_out = 8'hC5;
                    16'hF733: data_out = 8'hC4;
                    16'hF734: data_out = 8'hC3;
                    16'hF735: data_out = 8'hC2;
                    16'hF736: data_out = 8'hC1;
                    16'hF737: data_out = 8'hC0;
                    16'hF738: data_out = 8'hBF;
                    16'hF739: data_out = 8'hBE;
                    16'hF73A: data_out = 8'hBD;
                    16'hF73B: data_out = 8'hBC;
                    16'hF73C: data_out = 8'hBB;
                    16'hF73D: data_out = 8'hBA;
                    16'hF73E: data_out = 8'hB9;
                    16'hF73F: data_out = 8'hB8;
                    16'hF740: data_out = 8'hB7;
                    16'hF741: data_out = 8'hB6;
                    16'hF742: data_out = 8'hB5;
                    16'hF743: data_out = 8'hB4;
                    16'hF744: data_out = 8'hB3;
                    16'hF745: data_out = 8'hB2;
                    16'hF746: data_out = 8'hB1;
                    16'hF747: data_out = 8'hB0;
                    16'hF748: data_out = 8'hAF;
                    16'hF749: data_out = 8'hAE;
                    16'hF74A: data_out = 8'hAD;
                    16'hF74B: data_out = 8'hAC;
                    16'hF74C: data_out = 8'hAB;
                    16'hF74D: data_out = 8'hAA;
                    16'hF74E: data_out = 8'hA9;
                    16'hF74F: data_out = 8'hA8;
                    16'hF750: data_out = 8'hA7;
                    16'hF751: data_out = 8'hA6;
                    16'hF752: data_out = 8'hA5;
                    16'hF753: data_out = 8'hA4;
                    16'hF754: data_out = 8'hA3;
                    16'hF755: data_out = 8'hA2;
                    16'hF756: data_out = 8'hA1;
                    16'hF757: data_out = 8'hA0;
                    16'hF758: data_out = 8'h9F;
                    16'hF759: data_out = 8'h9E;
                    16'hF75A: data_out = 8'h9D;
                    16'hF75B: data_out = 8'h9C;
                    16'hF75C: data_out = 8'h9B;
                    16'hF75D: data_out = 8'h9A;
                    16'hF75E: data_out = 8'h99;
                    16'hF75F: data_out = 8'h98;
                    16'hF760: data_out = 8'h97;
                    16'hF761: data_out = 8'h96;
                    16'hF762: data_out = 8'h95;
                    16'hF763: data_out = 8'h94;
                    16'hF764: data_out = 8'h93;
                    16'hF765: data_out = 8'h92;
                    16'hF766: data_out = 8'h91;
                    16'hF767: data_out = 8'h90;
                    16'hF768: data_out = 8'h8F;
                    16'hF769: data_out = 8'h8E;
                    16'hF76A: data_out = 8'h8D;
                    16'hF76B: data_out = 8'h8C;
                    16'hF76C: data_out = 8'h8B;
                    16'hF76D: data_out = 8'h8A;
                    16'hF76E: data_out = 8'h89;
                    16'hF76F: data_out = 8'h88;
                    16'hF770: data_out = 8'h87;
                    16'hF771: data_out = 8'h86;
                    16'hF772: data_out = 8'h85;
                    16'hF773: data_out = 8'h84;
                    16'hF774: data_out = 8'h83;
                    16'hF775: data_out = 8'h82;
                    16'hF776: data_out = 8'h81;
                    16'hF777: data_out = 8'h0;
                    16'hF778: data_out = 8'h1;
                    16'hF779: data_out = 8'h2;
                    16'hF77A: data_out = 8'h3;
                    16'hF77B: data_out = 8'h4;
                    16'hF77C: data_out = 8'h5;
                    16'hF77D: data_out = 8'h6;
                    16'hF77E: data_out = 8'h7;
                    16'hF77F: data_out = 8'h8;
                    16'hF780: data_out = 8'hF7;
                    16'hF781: data_out = 8'hF8;
                    16'hF782: data_out = 8'hF9;
                    16'hF783: data_out = 8'hFA;
                    16'hF784: data_out = 8'hFB;
                    16'hF785: data_out = 8'hFC;
                    16'hF786: data_out = 8'hFD;
                    16'hF787: data_out = 8'hFE;
                    16'hF788: data_out = 8'hFF;
                    16'hF789: data_out = 8'h80;
                    16'hF78A: data_out = 8'h81;
                    16'hF78B: data_out = 8'h82;
                    16'hF78C: data_out = 8'h83;
                    16'hF78D: data_out = 8'h84;
                    16'hF78E: data_out = 8'h85;
                    16'hF78F: data_out = 8'h86;
                    16'hF790: data_out = 8'h87;
                    16'hF791: data_out = 8'h88;
                    16'hF792: data_out = 8'h89;
                    16'hF793: data_out = 8'h8A;
                    16'hF794: data_out = 8'h8B;
                    16'hF795: data_out = 8'h8C;
                    16'hF796: data_out = 8'h8D;
                    16'hF797: data_out = 8'h8E;
                    16'hF798: data_out = 8'h8F;
                    16'hF799: data_out = 8'h90;
                    16'hF79A: data_out = 8'h91;
                    16'hF79B: data_out = 8'h92;
                    16'hF79C: data_out = 8'h93;
                    16'hF79D: data_out = 8'h94;
                    16'hF79E: data_out = 8'h95;
                    16'hF79F: data_out = 8'h96;
                    16'hF7A0: data_out = 8'h97;
                    16'hF7A1: data_out = 8'h98;
                    16'hF7A2: data_out = 8'h99;
                    16'hF7A3: data_out = 8'h9A;
                    16'hF7A4: data_out = 8'h9B;
                    16'hF7A5: data_out = 8'h9C;
                    16'hF7A6: data_out = 8'h9D;
                    16'hF7A7: data_out = 8'h9E;
                    16'hF7A8: data_out = 8'h9F;
                    16'hF7A9: data_out = 8'hA0;
                    16'hF7AA: data_out = 8'hA1;
                    16'hF7AB: data_out = 8'hA2;
                    16'hF7AC: data_out = 8'hA3;
                    16'hF7AD: data_out = 8'hA4;
                    16'hF7AE: data_out = 8'hA5;
                    16'hF7AF: data_out = 8'hA6;
                    16'hF7B0: data_out = 8'hA7;
                    16'hF7B1: data_out = 8'hA8;
                    16'hF7B2: data_out = 8'hA9;
                    16'hF7B3: data_out = 8'hAA;
                    16'hF7B4: data_out = 8'hAB;
                    16'hF7B5: data_out = 8'hAC;
                    16'hF7B6: data_out = 8'hAD;
                    16'hF7B7: data_out = 8'hAE;
                    16'hF7B8: data_out = 8'hAF;
                    16'hF7B9: data_out = 8'hB0;
                    16'hF7BA: data_out = 8'hB1;
                    16'hF7BB: data_out = 8'hB2;
                    16'hF7BC: data_out = 8'hB3;
                    16'hF7BD: data_out = 8'hB4;
                    16'hF7BE: data_out = 8'hB5;
                    16'hF7BF: data_out = 8'hB6;
                    16'hF7C0: data_out = 8'hB7;
                    16'hF7C1: data_out = 8'hB8;
                    16'hF7C2: data_out = 8'hB9;
                    16'hF7C3: data_out = 8'hBA;
                    16'hF7C4: data_out = 8'hBB;
                    16'hF7C5: data_out = 8'hBC;
                    16'hF7C6: data_out = 8'hBD;
                    16'hF7C7: data_out = 8'hBE;
                    16'hF7C8: data_out = 8'hBF;
                    16'hF7C9: data_out = 8'hC0;
                    16'hF7CA: data_out = 8'hC1;
                    16'hF7CB: data_out = 8'hC2;
                    16'hF7CC: data_out = 8'hC3;
                    16'hF7CD: data_out = 8'hC4;
                    16'hF7CE: data_out = 8'hC5;
                    16'hF7CF: data_out = 8'hC6;
                    16'hF7D0: data_out = 8'hC7;
                    16'hF7D1: data_out = 8'hC8;
                    16'hF7D2: data_out = 8'hC9;
                    16'hF7D3: data_out = 8'hCA;
                    16'hF7D4: data_out = 8'hCB;
                    16'hF7D5: data_out = 8'hCC;
                    16'hF7D6: data_out = 8'hCD;
                    16'hF7D7: data_out = 8'hCE;
                    16'hF7D8: data_out = 8'hCF;
                    16'hF7D9: data_out = 8'hD0;
                    16'hF7DA: data_out = 8'hD1;
                    16'hF7DB: data_out = 8'hD2;
                    16'hF7DC: data_out = 8'hD3;
                    16'hF7DD: data_out = 8'hD4;
                    16'hF7DE: data_out = 8'hD5;
                    16'hF7DF: data_out = 8'hD6;
                    16'hF7E0: data_out = 8'hD7;
                    16'hF7E1: data_out = 8'hD8;
                    16'hF7E2: data_out = 8'hD9;
                    16'hF7E3: data_out = 8'hDA;
                    16'hF7E4: data_out = 8'hDB;
                    16'hF7E5: data_out = 8'hDC;
                    16'hF7E6: data_out = 8'hDD;
                    16'hF7E7: data_out = 8'hDE;
                    16'hF7E8: data_out = 8'hDF;
                    16'hF7E9: data_out = 8'hE0;
                    16'hF7EA: data_out = 8'hE1;
                    16'hF7EB: data_out = 8'hE2;
                    16'hF7EC: data_out = 8'hE3;
                    16'hF7ED: data_out = 8'hE4;
                    16'hF7EE: data_out = 8'hE5;
                    16'hF7EF: data_out = 8'hE6;
                    16'hF7F0: data_out = 8'hE7;
                    16'hF7F1: data_out = 8'hE8;
                    16'hF7F2: data_out = 8'hE9;
                    16'hF7F3: data_out = 8'hEA;
                    16'hF7F4: data_out = 8'hEB;
                    16'hF7F5: data_out = 8'hEC;
                    16'hF7F6: data_out = 8'hED;
                    16'hF7F7: data_out = 8'hEE;
                    16'hF7F8: data_out = 8'hEF;
                    16'hF7F9: data_out = 8'hF0;
                    16'hF7FA: data_out = 8'hF1;
                    16'hF7FB: data_out = 8'hF2;
                    16'hF7FC: data_out = 8'hF3;
                    16'hF7FD: data_out = 8'hF4;
                    16'hF7FE: data_out = 8'hF5;
                    16'hF7FF: data_out = 8'hF6;
                    16'hF800: data_out = 8'hF8;
                    16'hF801: data_out = 8'hF7;
                    16'hF802: data_out = 8'hF6;
                    16'hF803: data_out = 8'hF5;
                    16'hF804: data_out = 8'hF4;
                    16'hF805: data_out = 8'hF3;
                    16'hF806: data_out = 8'hF2;
                    16'hF807: data_out = 8'hF1;
                    16'hF808: data_out = 8'hF0;
                    16'hF809: data_out = 8'hEF;
                    16'hF80A: data_out = 8'hEE;
                    16'hF80B: data_out = 8'hED;
                    16'hF80C: data_out = 8'hEC;
                    16'hF80D: data_out = 8'hEB;
                    16'hF80E: data_out = 8'hEA;
                    16'hF80F: data_out = 8'hE9;
                    16'hF810: data_out = 8'hE8;
                    16'hF811: data_out = 8'hE7;
                    16'hF812: data_out = 8'hE6;
                    16'hF813: data_out = 8'hE5;
                    16'hF814: data_out = 8'hE4;
                    16'hF815: data_out = 8'hE3;
                    16'hF816: data_out = 8'hE2;
                    16'hF817: data_out = 8'hE1;
                    16'hF818: data_out = 8'hE0;
                    16'hF819: data_out = 8'hDF;
                    16'hF81A: data_out = 8'hDE;
                    16'hF81B: data_out = 8'hDD;
                    16'hF81C: data_out = 8'hDC;
                    16'hF81D: data_out = 8'hDB;
                    16'hF81E: data_out = 8'hDA;
                    16'hF81F: data_out = 8'hD9;
                    16'hF820: data_out = 8'hD8;
                    16'hF821: data_out = 8'hD7;
                    16'hF822: data_out = 8'hD6;
                    16'hF823: data_out = 8'hD5;
                    16'hF824: data_out = 8'hD4;
                    16'hF825: data_out = 8'hD3;
                    16'hF826: data_out = 8'hD2;
                    16'hF827: data_out = 8'hD1;
                    16'hF828: data_out = 8'hD0;
                    16'hF829: data_out = 8'hCF;
                    16'hF82A: data_out = 8'hCE;
                    16'hF82B: data_out = 8'hCD;
                    16'hF82C: data_out = 8'hCC;
                    16'hF82D: data_out = 8'hCB;
                    16'hF82E: data_out = 8'hCA;
                    16'hF82F: data_out = 8'hC9;
                    16'hF830: data_out = 8'hC8;
                    16'hF831: data_out = 8'hC7;
                    16'hF832: data_out = 8'hC6;
                    16'hF833: data_out = 8'hC5;
                    16'hF834: data_out = 8'hC4;
                    16'hF835: data_out = 8'hC3;
                    16'hF836: data_out = 8'hC2;
                    16'hF837: data_out = 8'hC1;
                    16'hF838: data_out = 8'hC0;
                    16'hF839: data_out = 8'hBF;
                    16'hF83A: data_out = 8'hBE;
                    16'hF83B: data_out = 8'hBD;
                    16'hF83C: data_out = 8'hBC;
                    16'hF83D: data_out = 8'hBB;
                    16'hF83E: data_out = 8'hBA;
                    16'hF83F: data_out = 8'hB9;
                    16'hF840: data_out = 8'hB8;
                    16'hF841: data_out = 8'hB7;
                    16'hF842: data_out = 8'hB6;
                    16'hF843: data_out = 8'hB5;
                    16'hF844: data_out = 8'hB4;
                    16'hF845: data_out = 8'hB3;
                    16'hF846: data_out = 8'hB2;
                    16'hF847: data_out = 8'hB1;
                    16'hF848: data_out = 8'hB0;
                    16'hF849: data_out = 8'hAF;
                    16'hF84A: data_out = 8'hAE;
                    16'hF84B: data_out = 8'hAD;
                    16'hF84C: data_out = 8'hAC;
                    16'hF84D: data_out = 8'hAB;
                    16'hF84E: data_out = 8'hAA;
                    16'hF84F: data_out = 8'hA9;
                    16'hF850: data_out = 8'hA8;
                    16'hF851: data_out = 8'hA7;
                    16'hF852: data_out = 8'hA6;
                    16'hF853: data_out = 8'hA5;
                    16'hF854: data_out = 8'hA4;
                    16'hF855: data_out = 8'hA3;
                    16'hF856: data_out = 8'hA2;
                    16'hF857: data_out = 8'hA1;
                    16'hF858: data_out = 8'hA0;
                    16'hF859: data_out = 8'h9F;
                    16'hF85A: data_out = 8'h9E;
                    16'hF85B: data_out = 8'h9D;
                    16'hF85C: data_out = 8'h9C;
                    16'hF85D: data_out = 8'h9B;
                    16'hF85E: data_out = 8'h9A;
                    16'hF85F: data_out = 8'h99;
                    16'hF860: data_out = 8'h98;
                    16'hF861: data_out = 8'h97;
                    16'hF862: data_out = 8'h96;
                    16'hF863: data_out = 8'h95;
                    16'hF864: data_out = 8'h94;
                    16'hF865: data_out = 8'h93;
                    16'hF866: data_out = 8'h92;
                    16'hF867: data_out = 8'h91;
                    16'hF868: data_out = 8'h90;
                    16'hF869: data_out = 8'h8F;
                    16'hF86A: data_out = 8'h8E;
                    16'hF86B: data_out = 8'h8D;
                    16'hF86C: data_out = 8'h8C;
                    16'hF86D: data_out = 8'h8B;
                    16'hF86E: data_out = 8'h8A;
                    16'hF86F: data_out = 8'h89;
                    16'hF870: data_out = 8'h88;
                    16'hF871: data_out = 8'h87;
                    16'hF872: data_out = 8'h86;
                    16'hF873: data_out = 8'h85;
                    16'hF874: data_out = 8'h84;
                    16'hF875: data_out = 8'h83;
                    16'hF876: data_out = 8'h82;
                    16'hF877: data_out = 8'h81;
                    16'hF878: data_out = 8'h0;
                    16'hF879: data_out = 8'h1;
                    16'hF87A: data_out = 8'h2;
                    16'hF87B: data_out = 8'h3;
                    16'hF87C: data_out = 8'h4;
                    16'hF87D: data_out = 8'h5;
                    16'hF87E: data_out = 8'h6;
                    16'hF87F: data_out = 8'h7;
                    16'hF880: data_out = 8'hF8;
                    16'hF881: data_out = 8'hF9;
                    16'hF882: data_out = 8'hFA;
                    16'hF883: data_out = 8'hFB;
                    16'hF884: data_out = 8'hFC;
                    16'hF885: data_out = 8'hFD;
                    16'hF886: data_out = 8'hFE;
                    16'hF887: data_out = 8'hFF;
                    16'hF888: data_out = 8'h80;
                    16'hF889: data_out = 8'h81;
                    16'hF88A: data_out = 8'h82;
                    16'hF88B: data_out = 8'h83;
                    16'hF88C: data_out = 8'h84;
                    16'hF88D: data_out = 8'h85;
                    16'hF88E: data_out = 8'h86;
                    16'hF88F: data_out = 8'h87;
                    16'hF890: data_out = 8'h88;
                    16'hF891: data_out = 8'h89;
                    16'hF892: data_out = 8'h8A;
                    16'hF893: data_out = 8'h8B;
                    16'hF894: data_out = 8'h8C;
                    16'hF895: data_out = 8'h8D;
                    16'hF896: data_out = 8'h8E;
                    16'hF897: data_out = 8'h8F;
                    16'hF898: data_out = 8'h90;
                    16'hF899: data_out = 8'h91;
                    16'hF89A: data_out = 8'h92;
                    16'hF89B: data_out = 8'h93;
                    16'hF89C: data_out = 8'h94;
                    16'hF89D: data_out = 8'h95;
                    16'hF89E: data_out = 8'h96;
                    16'hF89F: data_out = 8'h97;
                    16'hF8A0: data_out = 8'h98;
                    16'hF8A1: data_out = 8'h99;
                    16'hF8A2: data_out = 8'h9A;
                    16'hF8A3: data_out = 8'h9B;
                    16'hF8A4: data_out = 8'h9C;
                    16'hF8A5: data_out = 8'h9D;
                    16'hF8A6: data_out = 8'h9E;
                    16'hF8A7: data_out = 8'h9F;
                    16'hF8A8: data_out = 8'hA0;
                    16'hF8A9: data_out = 8'hA1;
                    16'hF8AA: data_out = 8'hA2;
                    16'hF8AB: data_out = 8'hA3;
                    16'hF8AC: data_out = 8'hA4;
                    16'hF8AD: data_out = 8'hA5;
                    16'hF8AE: data_out = 8'hA6;
                    16'hF8AF: data_out = 8'hA7;
                    16'hF8B0: data_out = 8'hA8;
                    16'hF8B1: data_out = 8'hA9;
                    16'hF8B2: data_out = 8'hAA;
                    16'hF8B3: data_out = 8'hAB;
                    16'hF8B4: data_out = 8'hAC;
                    16'hF8B5: data_out = 8'hAD;
                    16'hF8B6: data_out = 8'hAE;
                    16'hF8B7: data_out = 8'hAF;
                    16'hF8B8: data_out = 8'hB0;
                    16'hF8B9: data_out = 8'hB1;
                    16'hF8BA: data_out = 8'hB2;
                    16'hF8BB: data_out = 8'hB3;
                    16'hF8BC: data_out = 8'hB4;
                    16'hF8BD: data_out = 8'hB5;
                    16'hF8BE: data_out = 8'hB6;
                    16'hF8BF: data_out = 8'hB7;
                    16'hF8C0: data_out = 8'hB8;
                    16'hF8C1: data_out = 8'hB9;
                    16'hF8C2: data_out = 8'hBA;
                    16'hF8C3: data_out = 8'hBB;
                    16'hF8C4: data_out = 8'hBC;
                    16'hF8C5: data_out = 8'hBD;
                    16'hF8C6: data_out = 8'hBE;
                    16'hF8C7: data_out = 8'hBF;
                    16'hF8C8: data_out = 8'hC0;
                    16'hF8C9: data_out = 8'hC1;
                    16'hF8CA: data_out = 8'hC2;
                    16'hF8CB: data_out = 8'hC3;
                    16'hF8CC: data_out = 8'hC4;
                    16'hF8CD: data_out = 8'hC5;
                    16'hF8CE: data_out = 8'hC6;
                    16'hF8CF: data_out = 8'hC7;
                    16'hF8D0: data_out = 8'hC8;
                    16'hF8D1: data_out = 8'hC9;
                    16'hF8D2: data_out = 8'hCA;
                    16'hF8D3: data_out = 8'hCB;
                    16'hF8D4: data_out = 8'hCC;
                    16'hF8D5: data_out = 8'hCD;
                    16'hF8D6: data_out = 8'hCE;
                    16'hF8D7: data_out = 8'hCF;
                    16'hF8D8: data_out = 8'hD0;
                    16'hF8D9: data_out = 8'hD1;
                    16'hF8DA: data_out = 8'hD2;
                    16'hF8DB: data_out = 8'hD3;
                    16'hF8DC: data_out = 8'hD4;
                    16'hF8DD: data_out = 8'hD5;
                    16'hF8DE: data_out = 8'hD6;
                    16'hF8DF: data_out = 8'hD7;
                    16'hF8E0: data_out = 8'hD8;
                    16'hF8E1: data_out = 8'hD9;
                    16'hF8E2: data_out = 8'hDA;
                    16'hF8E3: data_out = 8'hDB;
                    16'hF8E4: data_out = 8'hDC;
                    16'hF8E5: data_out = 8'hDD;
                    16'hF8E6: data_out = 8'hDE;
                    16'hF8E7: data_out = 8'hDF;
                    16'hF8E8: data_out = 8'hE0;
                    16'hF8E9: data_out = 8'hE1;
                    16'hF8EA: data_out = 8'hE2;
                    16'hF8EB: data_out = 8'hE3;
                    16'hF8EC: data_out = 8'hE4;
                    16'hF8ED: data_out = 8'hE5;
                    16'hF8EE: data_out = 8'hE6;
                    16'hF8EF: data_out = 8'hE7;
                    16'hF8F0: data_out = 8'hE8;
                    16'hF8F1: data_out = 8'hE9;
                    16'hF8F2: data_out = 8'hEA;
                    16'hF8F3: data_out = 8'hEB;
                    16'hF8F4: data_out = 8'hEC;
                    16'hF8F5: data_out = 8'hED;
                    16'hF8F6: data_out = 8'hEE;
                    16'hF8F7: data_out = 8'hEF;
                    16'hF8F8: data_out = 8'hF0;
                    16'hF8F9: data_out = 8'hF1;
                    16'hF8FA: data_out = 8'hF2;
                    16'hF8FB: data_out = 8'hF3;
                    16'hF8FC: data_out = 8'hF4;
                    16'hF8FD: data_out = 8'hF5;
                    16'hF8FE: data_out = 8'hF6;
                    16'hF8FF: data_out = 8'hF7;
                    16'hF900: data_out = 8'hF9;
                    16'hF901: data_out = 8'hF8;
                    16'hF902: data_out = 8'hF7;
                    16'hF903: data_out = 8'hF6;
                    16'hF904: data_out = 8'hF5;
                    16'hF905: data_out = 8'hF4;
                    16'hF906: data_out = 8'hF3;
                    16'hF907: data_out = 8'hF2;
                    16'hF908: data_out = 8'hF1;
                    16'hF909: data_out = 8'hF0;
                    16'hF90A: data_out = 8'hEF;
                    16'hF90B: data_out = 8'hEE;
                    16'hF90C: data_out = 8'hED;
                    16'hF90D: data_out = 8'hEC;
                    16'hF90E: data_out = 8'hEB;
                    16'hF90F: data_out = 8'hEA;
                    16'hF910: data_out = 8'hE9;
                    16'hF911: data_out = 8'hE8;
                    16'hF912: data_out = 8'hE7;
                    16'hF913: data_out = 8'hE6;
                    16'hF914: data_out = 8'hE5;
                    16'hF915: data_out = 8'hE4;
                    16'hF916: data_out = 8'hE3;
                    16'hF917: data_out = 8'hE2;
                    16'hF918: data_out = 8'hE1;
                    16'hF919: data_out = 8'hE0;
                    16'hF91A: data_out = 8'hDF;
                    16'hF91B: data_out = 8'hDE;
                    16'hF91C: data_out = 8'hDD;
                    16'hF91D: data_out = 8'hDC;
                    16'hF91E: data_out = 8'hDB;
                    16'hF91F: data_out = 8'hDA;
                    16'hF920: data_out = 8'hD9;
                    16'hF921: data_out = 8'hD8;
                    16'hF922: data_out = 8'hD7;
                    16'hF923: data_out = 8'hD6;
                    16'hF924: data_out = 8'hD5;
                    16'hF925: data_out = 8'hD4;
                    16'hF926: data_out = 8'hD3;
                    16'hF927: data_out = 8'hD2;
                    16'hF928: data_out = 8'hD1;
                    16'hF929: data_out = 8'hD0;
                    16'hF92A: data_out = 8'hCF;
                    16'hF92B: data_out = 8'hCE;
                    16'hF92C: data_out = 8'hCD;
                    16'hF92D: data_out = 8'hCC;
                    16'hF92E: data_out = 8'hCB;
                    16'hF92F: data_out = 8'hCA;
                    16'hF930: data_out = 8'hC9;
                    16'hF931: data_out = 8'hC8;
                    16'hF932: data_out = 8'hC7;
                    16'hF933: data_out = 8'hC6;
                    16'hF934: data_out = 8'hC5;
                    16'hF935: data_out = 8'hC4;
                    16'hF936: data_out = 8'hC3;
                    16'hF937: data_out = 8'hC2;
                    16'hF938: data_out = 8'hC1;
                    16'hF939: data_out = 8'hC0;
                    16'hF93A: data_out = 8'hBF;
                    16'hF93B: data_out = 8'hBE;
                    16'hF93C: data_out = 8'hBD;
                    16'hF93D: data_out = 8'hBC;
                    16'hF93E: data_out = 8'hBB;
                    16'hF93F: data_out = 8'hBA;
                    16'hF940: data_out = 8'hB9;
                    16'hF941: data_out = 8'hB8;
                    16'hF942: data_out = 8'hB7;
                    16'hF943: data_out = 8'hB6;
                    16'hF944: data_out = 8'hB5;
                    16'hF945: data_out = 8'hB4;
                    16'hF946: data_out = 8'hB3;
                    16'hF947: data_out = 8'hB2;
                    16'hF948: data_out = 8'hB1;
                    16'hF949: data_out = 8'hB0;
                    16'hF94A: data_out = 8'hAF;
                    16'hF94B: data_out = 8'hAE;
                    16'hF94C: data_out = 8'hAD;
                    16'hF94D: data_out = 8'hAC;
                    16'hF94E: data_out = 8'hAB;
                    16'hF94F: data_out = 8'hAA;
                    16'hF950: data_out = 8'hA9;
                    16'hF951: data_out = 8'hA8;
                    16'hF952: data_out = 8'hA7;
                    16'hF953: data_out = 8'hA6;
                    16'hF954: data_out = 8'hA5;
                    16'hF955: data_out = 8'hA4;
                    16'hF956: data_out = 8'hA3;
                    16'hF957: data_out = 8'hA2;
                    16'hF958: data_out = 8'hA1;
                    16'hF959: data_out = 8'hA0;
                    16'hF95A: data_out = 8'h9F;
                    16'hF95B: data_out = 8'h9E;
                    16'hF95C: data_out = 8'h9D;
                    16'hF95D: data_out = 8'h9C;
                    16'hF95E: data_out = 8'h9B;
                    16'hF95F: data_out = 8'h9A;
                    16'hF960: data_out = 8'h99;
                    16'hF961: data_out = 8'h98;
                    16'hF962: data_out = 8'h97;
                    16'hF963: data_out = 8'h96;
                    16'hF964: data_out = 8'h95;
                    16'hF965: data_out = 8'h94;
                    16'hF966: data_out = 8'h93;
                    16'hF967: data_out = 8'h92;
                    16'hF968: data_out = 8'h91;
                    16'hF969: data_out = 8'h90;
                    16'hF96A: data_out = 8'h8F;
                    16'hF96B: data_out = 8'h8E;
                    16'hF96C: data_out = 8'h8D;
                    16'hF96D: data_out = 8'h8C;
                    16'hF96E: data_out = 8'h8B;
                    16'hF96F: data_out = 8'h8A;
                    16'hF970: data_out = 8'h89;
                    16'hF971: data_out = 8'h88;
                    16'hF972: data_out = 8'h87;
                    16'hF973: data_out = 8'h86;
                    16'hF974: data_out = 8'h85;
                    16'hF975: data_out = 8'h84;
                    16'hF976: data_out = 8'h83;
                    16'hF977: data_out = 8'h82;
                    16'hF978: data_out = 8'h81;
                    16'hF979: data_out = 8'h0;
                    16'hF97A: data_out = 8'h1;
                    16'hF97B: data_out = 8'h2;
                    16'hF97C: data_out = 8'h3;
                    16'hF97D: data_out = 8'h4;
                    16'hF97E: data_out = 8'h5;
                    16'hF97F: data_out = 8'h6;
                    16'hF980: data_out = 8'hF9;
                    16'hF981: data_out = 8'hFA;
                    16'hF982: data_out = 8'hFB;
                    16'hF983: data_out = 8'hFC;
                    16'hF984: data_out = 8'hFD;
                    16'hF985: data_out = 8'hFE;
                    16'hF986: data_out = 8'hFF;
                    16'hF987: data_out = 8'h80;
                    16'hF988: data_out = 8'h81;
                    16'hF989: data_out = 8'h82;
                    16'hF98A: data_out = 8'h83;
                    16'hF98B: data_out = 8'h84;
                    16'hF98C: data_out = 8'h85;
                    16'hF98D: data_out = 8'h86;
                    16'hF98E: data_out = 8'h87;
                    16'hF98F: data_out = 8'h88;
                    16'hF990: data_out = 8'h89;
                    16'hF991: data_out = 8'h8A;
                    16'hF992: data_out = 8'h8B;
                    16'hF993: data_out = 8'h8C;
                    16'hF994: data_out = 8'h8D;
                    16'hF995: data_out = 8'h8E;
                    16'hF996: data_out = 8'h8F;
                    16'hF997: data_out = 8'h90;
                    16'hF998: data_out = 8'h91;
                    16'hF999: data_out = 8'h92;
                    16'hF99A: data_out = 8'h93;
                    16'hF99B: data_out = 8'h94;
                    16'hF99C: data_out = 8'h95;
                    16'hF99D: data_out = 8'h96;
                    16'hF99E: data_out = 8'h97;
                    16'hF99F: data_out = 8'h98;
                    16'hF9A0: data_out = 8'h99;
                    16'hF9A1: data_out = 8'h9A;
                    16'hF9A2: data_out = 8'h9B;
                    16'hF9A3: data_out = 8'h9C;
                    16'hF9A4: data_out = 8'h9D;
                    16'hF9A5: data_out = 8'h9E;
                    16'hF9A6: data_out = 8'h9F;
                    16'hF9A7: data_out = 8'hA0;
                    16'hF9A8: data_out = 8'hA1;
                    16'hF9A9: data_out = 8'hA2;
                    16'hF9AA: data_out = 8'hA3;
                    16'hF9AB: data_out = 8'hA4;
                    16'hF9AC: data_out = 8'hA5;
                    16'hF9AD: data_out = 8'hA6;
                    16'hF9AE: data_out = 8'hA7;
                    16'hF9AF: data_out = 8'hA8;
                    16'hF9B0: data_out = 8'hA9;
                    16'hF9B1: data_out = 8'hAA;
                    16'hF9B2: data_out = 8'hAB;
                    16'hF9B3: data_out = 8'hAC;
                    16'hF9B4: data_out = 8'hAD;
                    16'hF9B5: data_out = 8'hAE;
                    16'hF9B6: data_out = 8'hAF;
                    16'hF9B7: data_out = 8'hB0;
                    16'hF9B8: data_out = 8'hB1;
                    16'hF9B9: data_out = 8'hB2;
                    16'hF9BA: data_out = 8'hB3;
                    16'hF9BB: data_out = 8'hB4;
                    16'hF9BC: data_out = 8'hB5;
                    16'hF9BD: data_out = 8'hB6;
                    16'hF9BE: data_out = 8'hB7;
                    16'hF9BF: data_out = 8'hB8;
                    16'hF9C0: data_out = 8'hB9;
                    16'hF9C1: data_out = 8'hBA;
                    16'hF9C2: data_out = 8'hBB;
                    16'hF9C3: data_out = 8'hBC;
                    16'hF9C4: data_out = 8'hBD;
                    16'hF9C5: data_out = 8'hBE;
                    16'hF9C6: data_out = 8'hBF;
                    16'hF9C7: data_out = 8'hC0;
                    16'hF9C8: data_out = 8'hC1;
                    16'hF9C9: data_out = 8'hC2;
                    16'hF9CA: data_out = 8'hC3;
                    16'hF9CB: data_out = 8'hC4;
                    16'hF9CC: data_out = 8'hC5;
                    16'hF9CD: data_out = 8'hC6;
                    16'hF9CE: data_out = 8'hC7;
                    16'hF9CF: data_out = 8'hC8;
                    16'hF9D0: data_out = 8'hC9;
                    16'hF9D1: data_out = 8'hCA;
                    16'hF9D2: data_out = 8'hCB;
                    16'hF9D3: data_out = 8'hCC;
                    16'hF9D4: data_out = 8'hCD;
                    16'hF9D5: data_out = 8'hCE;
                    16'hF9D6: data_out = 8'hCF;
                    16'hF9D7: data_out = 8'hD0;
                    16'hF9D8: data_out = 8'hD1;
                    16'hF9D9: data_out = 8'hD2;
                    16'hF9DA: data_out = 8'hD3;
                    16'hF9DB: data_out = 8'hD4;
                    16'hF9DC: data_out = 8'hD5;
                    16'hF9DD: data_out = 8'hD6;
                    16'hF9DE: data_out = 8'hD7;
                    16'hF9DF: data_out = 8'hD8;
                    16'hF9E0: data_out = 8'hD9;
                    16'hF9E1: data_out = 8'hDA;
                    16'hF9E2: data_out = 8'hDB;
                    16'hF9E3: data_out = 8'hDC;
                    16'hF9E4: data_out = 8'hDD;
                    16'hF9E5: data_out = 8'hDE;
                    16'hF9E6: data_out = 8'hDF;
                    16'hF9E7: data_out = 8'hE0;
                    16'hF9E8: data_out = 8'hE1;
                    16'hF9E9: data_out = 8'hE2;
                    16'hF9EA: data_out = 8'hE3;
                    16'hF9EB: data_out = 8'hE4;
                    16'hF9EC: data_out = 8'hE5;
                    16'hF9ED: data_out = 8'hE6;
                    16'hF9EE: data_out = 8'hE7;
                    16'hF9EF: data_out = 8'hE8;
                    16'hF9F0: data_out = 8'hE9;
                    16'hF9F1: data_out = 8'hEA;
                    16'hF9F2: data_out = 8'hEB;
                    16'hF9F3: data_out = 8'hEC;
                    16'hF9F4: data_out = 8'hED;
                    16'hF9F5: data_out = 8'hEE;
                    16'hF9F6: data_out = 8'hEF;
                    16'hF9F7: data_out = 8'hF0;
                    16'hF9F8: data_out = 8'hF1;
                    16'hF9F9: data_out = 8'hF2;
                    16'hF9FA: data_out = 8'hF3;
                    16'hF9FB: data_out = 8'hF4;
                    16'hF9FC: data_out = 8'hF5;
                    16'hF9FD: data_out = 8'hF6;
                    16'hF9FE: data_out = 8'hF7;
                    16'hF9FF: data_out = 8'hF8;
                    16'hFA00: data_out = 8'hFA;
                    16'hFA01: data_out = 8'hF9;
                    16'hFA02: data_out = 8'hF8;
                    16'hFA03: data_out = 8'hF7;
                    16'hFA04: data_out = 8'hF6;
                    16'hFA05: data_out = 8'hF5;
                    16'hFA06: data_out = 8'hF4;
                    16'hFA07: data_out = 8'hF3;
                    16'hFA08: data_out = 8'hF2;
                    16'hFA09: data_out = 8'hF1;
                    16'hFA0A: data_out = 8'hF0;
                    16'hFA0B: data_out = 8'hEF;
                    16'hFA0C: data_out = 8'hEE;
                    16'hFA0D: data_out = 8'hED;
                    16'hFA0E: data_out = 8'hEC;
                    16'hFA0F: data_out = 8'hEB;
                    16'hFA10: data_out = 8'hEA;
                    16'hFA11: data_out = 8'hE9;
                    16'hFA12: data_out = 8'hE8;
                    16'hFA13: data_out = 8'hE7;
                    16'hFA14: data_out = 8'hE6;
                    16'hFA15: data_out = 8'hE5;
                    16'hFA16: data_out = 8'hE4;
                    16'hFA17: data_out = 8'hE3;
                    16'hFA18: data_out = 8'hE2;
                    16'hFA19: data_out = 8'hE1;
                    16'hFA1A: data_out = 8'hE0;
                    16'hFA1B: data_out = 8'hDF;
                    16'hFA1C: data_out = 8'hDE;
                    16'hFA1D: data_out = 8'hDD;
                    16'hFA1E: data_out = 8'hDC;
                    16'hFA1F: data_out = 8'hDB;
                    16'hFA20: data_out = 8'hDA;
                    16'hFA21: data_out = 8'hD9;
                    16'hFA22: data_out = 8'hD8;
                    16'hFA23: data_out = 8'hD7;
                    16'hFA24: data_out = 8'hD6;
                    16'hFA25: data_out = 8'hD5;
                    16'hFA26: data_out = 8'hD4;
                    16'hFA27: data_out = 8'hD3;
                    16'hFA28: data_out = 8'hD2;
                    16'hFA29: data_out = 8'hD1;
                    16'hFA2A: data_out = 8'hD0;
                    16'hFA2B: data_out = 8'hCF;
                    16'hFA2C: data_out = 8'hCE;
                    16'hFA2D: data_out = 8'hCD;
                    16'hFA2E: data_out = 8'hCC;
                    16'hFA2F: data_out = 8'hCB;
                    16'hFA30: data_out = 8'hCA;
                    16'hFA31: data_out = 8'hC9;
                    16'hFA32: data_out = 8'hC8;
                    16'hFA33: data_out = 8'hC7;
                    16'hFA34: data_out = 8'hC6;
                    16'hFA35: data_out = 8'hC5;
                    16'hFA36: data_out = 8'hC4;
                    16'hFA37: data_out = 8'hC3;
                    16'hFA38: data_out = 8'hC2;
                    16'hFA39: data_out = 8'hC1;
                    16'hFA3A: data_out = 8'hC0;
                    16'hFA3B: data_out = 8'hBF;
                    16'hFA3C: data_out = 8'hBE;
                    16'hFA3D: data_out = 8'hBD;
                    16'hFA3E: data_out = 8'hBC;
                    16'hFA3F: data_out = 8'hBB;
                    16'hFA40: data_out = 8'hBA;
                    16'hFA41: data_out = 8'hB9;
                    16'hFA42: data_out = 8'hB8;
                    16'hFA43: data_out = 8'hB7;
                    16'hFA44: data_out = 8'hB6;
                    16'hFA45: data_out = 8'hB5;
                    16'hFA46: data_out = 8'hB4;
                    16'hFA47: data_out = 8'hB3;
                    16'hFA48: data_out = 8'hB2;
                    16'hFA49: data_out = 8'hB1;
                    16'hFA4A: data_out = 8'hB0;
                    16'hFA4B: data_out = 8'hAF;
                    16'hFA4C: data_out = 8'hAE;
                    16'hFA4D: data_out = 8'hAD;
                    16'hFA4E: data_out = 8'hAC;
                    16'hFA4F: data_out = 8'hAB;
                    16'hFA50: data_out = 8'hAA;
                    16'hFA51: data_out = 8'hA9;
                    16'hFA52: data_out = 8'hA8;
                    16'hFA53: data_out = 8'hA7;
                    16'hFA54: data_out = 8'hA6;
                    16'hFA55: data_out = 8'hA5;
                    16'hFA56: data_out = 8'hA4;
                    16'hFA57: data_out = 8'hA3;
                    16'hFA58: data_out = 8'hA2;
                    16'hFA59: data_out = 8'hA1;
                    16'hFA5A: data_out = 8'hA0;
                    16'hFA5B: data_out = 8'h9F;
                    16'hFA5C: data_out = 8'h9E;
                    16'hFA5D: data_out = 8'h9D;
                    16'hFA5E: data_out = 8'h9C;
                    16'hFA5F: data_out = 8'h9B;
                    16'hFA60: data_out = 8'h9A;
                    16'hFA61: data_out = 8'h99;
                    16'hFA62: data_out = 8'h98;
                    16'hFA63: data_out = 8'h97;
                    16'hFA64: data_out = 8'h96;
                    16'hFA65: data_out = 8'h95;
                    16'hFA66: data_out = 8'h94;
                    16'hFA67: data_out = 8'h93;
                    16'hFA68: data_out = 8'h92;
                    16'hFA69: data_out = 8'h91;
                    16'hFA6A: data_out = 8'h90;
                    16'hFA6B: data_out = 8'h8F;
                    16'hFA6C: data_out = 8'h8E;
                    16'hFA6D: data_out = 8'h8D;
                    16'hFA6E: data_out = 8'h8C;
                    16'hFA6F: data_out = 8'h8B;
                    16'hFA70: data_out = 8'h8A;
                    16'hFA71: data_out = 8'h89;
                    16'hFA72: data_out = 8'h88;
                    16'hFA73: data_out = 8'h87;
                    16'hFA74: data_out = 8'h86;
                    16'hFA75: data_out = 8'h85;
                    16'hFA76: data_out = 8'h84;
                    16'hFA77: data_out = 8'h83;
                    16'hFA78: data_out = 8'h82;
                    16'hFA79: data_out = 8'h81;
                    16'hFA7A: data_out = 8'h0;
                    16'hFA7B: data_out = 8'h1;
                    16'hFA7C: data_out = 8'h2;
                    16'hFA7D: data_out = 8'h3;
                    16'hFA7E: data_out = 8'h4;
                    16'hFA7F: data_out = 8'h5;
                    16'hFA80: data_out = 8'hFA;
                    16'hFA81: data_out = 8'hFB;
                    16'hFA82: data_out = 8'hFC;
                    16'hFA83: data_out = 8'hFD;
                    16'hFA84: data_out = 8'hFE;
                    16'hFA85: data_out = 8'hFF;
                    16'hFA86: data_out = 8'h80;
                    16'hFA87: data_out = 8'h81;
                    16'hFA88: data_out = 8'h82;
                    16'hFA89: data_out = 8'h83;
                    16'hFA8A: data_out = 8'h84;
                    16'hFA8B: data_out = 8'h85;
                    16'hFA8C: data_out = 8'h86;
                    16'hFA8D: data_out = 8'h87;
                    16'hFA8E: data_out = 8'h88;
                    16'hFA8F: data_out = 8'h89;
                    16'hFA90: data_out = 8'h8A;
                    16'hFA91: data_out = 8'h8B;
                    16'hFA92: data_out = 8'h8C;
                    16'hFA93: data_out = 8'h8D;
                    16'hFA94: data_out = 8'h8E;
                    16'hFA95: data_out = 8'h8F;
                    16'hFA96: data_out = 8'h90;
                    16'hFA97: data_out = 8'h91;
                    16'hFA98: data_out = 8'h92;
                    16'hFA99: data_out = 8'h93;
                    16'hFA9A: data_out = 8'h94;
                    16'hFA9B: data_out = 8'h95;
                    16'hFA9C: data_out = 8'h96;
                    16'hFA9D: data_out = 8'h97;
                    16'hFA9E: data_out = 8'h98;
                    16'hFA9F: data_out = 8'h99;
                    16'hFAA0: data_out = 8'h9A;
                    16'hFAA1: data_out = 8'h9B;
                    16'hFAA2: data_out = 8'h9C;
                    16'hFAA3: data_out = 8'h9D;
                    16'hFAA4: data_out = 8'h9E;
                    16'hFAA5: data_out = 8'h9F;
                    16'hFAA6: data_out = 8'hA0;
                    16'hFAA7: data_out = 8'hA1;
                    16'hFAA8: data_out = 8'hA2;
                    16'hFAA9: data_out = 8'hA3;
                    16'hFAAA: data_out = 8'hA4;
                    16'hFAAB: data_out = 8'hA5;
                    16'hFAAC: data_out = 8'hA6;
                    16'hFAAD: data_out = 8'hA7;
                    16'hFAAE: data_out = 8'hA8;
                    16'hFAAF: data_out = 8'hA9;
                    16'hFAB0: data_out = 8'hAA;
                    16'hFAB1: data_out = 8'hAB;
                    16'hFAB2: data_out = 8'hAC;
                    16'hFAB3: data_out = 8'hAD;
                    16'hFAB4: data_out = 8'hAE;
                    16'hFAB5: data_out = 8'hAF;
                    16'hFAB6: data_out = 8'hB0;
                    16'hFAB7: data_out = 8'hB1;
                    16'hFAB8: data_out = 8'hB2;
                    16'hFAB9: data_out = 8'hB3;
                    16'hFABA: data_out = 8'hB4;
                    16'hFABB: data_out = 8'hB5;
                    16'hFABC: data_out = 8'hB6;
                    16'hFABD: data_out = 8'hB7;
                    16'hFABE: data_out = 8'hB8;
                    16'hFABF: data_out = 8'hB9;
                    16'hFAC0: data_out = 8'hBA;
                    16'hFAC1: data_out = 8'hBB;
                    16'hFAC2: data_out = 8'hBC;
                    16'hFAC3: data_out = 8'hBD;
                    16'hFAC4: data_out = 8'hBE;
                    16'hFAC5: data_out = 8'hBF;
                    16'hFAC6: data_out = 8'hC0;
                    16'hFAC7: data_out = 8'hC1;
                    16'hFAC8: data_out = 8'hC2;
                    16'hFAC9: data_out = 8'hC3;
                    16'hFACA: data_out = 8'hC4;
                    16'hFACB: data_out = 8'hC5;
                    16'hFACC: data_out = 8'hC6;
                    16'hFACD: data_out = 8'hC7;
                    16'hFACE: data_out = 8'hC8;
                    16'hFACF: data_out = 8'hC9;
                    16'hFAD0: data_out = 8'hCA;
                    16'hFAD1: data_out = 8'hCB;
                    16'hFAD2: data_out = 8'hCC;
                    16'hFAD3: data_out = 8'hCD;
                    16'hFAD4: data_out = 8'hCE;
                    16'hFAD5: data_out = 8'hCF;
                    16'hFAD6: data_out = 8'hD0;
                    16'hFAD7: data_out = 8'hD1;
                    16'hFAD8: data_out = 8'hD2;
                    16'hFAD9: data_out = 8'hD3;
                    16'hFADA: data_out = 8'hD4;
                    16'hFADB: data_out = 8'hD5;
                    16'hFADC: data_out = 8'hD6;
                    16'hFADD: data_out = 8'hD7;
                    16'hFADE: data_out = 8'hD8;
                    16'hFADF: data_out = 8'hD9;
                    16'hFAE0: data_out = 8'hDA;
                    16'hFAE1: data_out = 8'hDB;
                    16'hFAE2: data_out = 8'hDC;
                    16'hFAE3: data_out = 8'hDD;
                    16'hFAE4: data_out = 8'hDE;
                    16'hFAE5: data_out = 8'hDF;
                    16'hFAE6: data_out = 8'hE0;
                    16'hFAE7: data_out = 8'hE1;
                    16'hFAE8: data_out = 8'hE2;
                    16'hFAE9: data_out = 8'hE3;
                    16'hFAEA: data_out = 8'hE4;
                    16'hFAEB: data_out = 8'hE5;
                    16'hFAEC: data_out = 8'hE6;
                    16'hFAED: data_out = 8'hE7;
                    16'hFAEE: data_out = 8'hE8;
                    16'hFAEF: data_out = 8'hE9;
                    16'hFAF0: data_out = 8'hEA;
                    16'hFAF1: data_out = 8'hEB;
                    16'hFAF2: data_out = 8'hEC;
                    16'hFAF3: data_out = 8'hED;
                    16'hFAF4: data_out = 8'hEE;
                    16'hFAF5: data_out = 8'hEF;
                    16'hFAF6: data_out = 8'hF0;
                    16'hFAF7: data_out = 8'hF1;
                    16'hFAF8: data_out = 8'hF2;
                    16'hFAF9: data_out = 8'hF3;
                    16'hFAFA: data_out = 8'hF4;
                    16'hFAFB: data_out = 8'hF5;
                    16'hFAFC: data_out = 8'hF6;
                    16'hFAFD: data_out = 8'hF7;
                    16'hFAFE: data_out = 8'hF8;
                    16'hFAFF: data_out = 8'hF9;
                    16'hFB00: data_out = 8'hFB;
                    16'hFB01: data_out = 8'hFA;
                    16'hFB02: data_out = 8'hF9;
                    16'hFB03: data_out = 8'hF8;
                    16'hFB04: data_out = 8'hF7;
                    16'hFB05: data_out = 8'hF6;
                    16'hFB06: data_out = 8'hF5;
                    16'hFB07: data_out = 8'hF4;
                    16'hFB08: data_out = 8'hF3;
                    16'hFB09: data_out = 8'hF2;
                    16'hFB0A: data_out = 8'hF1;
                    16'hFB0B: data_out = 8'hF0;
                    16'hFB0C: data_out = 8'hEF;
                    16'hFB0D: data_out = 8'hEE;
                    16'hFB0E: data_out = 8'hED;
                    16'hFB0F: data_out = 8'hEC;
                    16'hFB10: data_out = 8'hEB;
                    16'hFB11: data_out = 8'hEA;
                    16'hFB12: data_out = 8'hE9;
                    16'hFB13: data_out = 8'hE8;
                    16'hFB14: data_out = 8'hE7;
                    16'hFB15: data_out = 8'hE6;
                    16'hFB16: data_out = 8'hE5;
                    16'hFB17: data_out = 8'hE4;
                    16'hFB18: data_out = 8'hE3;
                    16'hFB19: data_out = 8'hE2;
                    16'hFB1A: data_out = 8'hE1;
                    16'hFB1B: data_out = 8'hE0;
                    16'hFB1C: data_out = 8'hDF;
                    16'hFB1D: data_out = 8'hDE;
                    16'hFB1E: data_out = 8'hDD;
                    16'hFB1F: data_out = 8'hDC;
                    16'hFB20: data_out = 8'hDB;
                    16'hFB21: data_out = 8'hDA;
                    16'hFB22: data_out = 8'hD9;
                    16'hFB23: data_out = 8'hD8;
                    16'hFB24: data_out = 8'hD7;
                    16'hFB25: data_out = 8'hD6;
                    16'hFB26: data_out = 8'hD5;
                    16'hFB27: data_out = 8'hD4;
                    16'hFB28: data_out = 8'hD3;
                    16'hFB29: data_out = 8'hD2;
                    16'hFB2A: data_out = 8'hD1;
                    16'hFB2B: data_out = 8'hD0;
                    16'hFB2C: data_out = 8'hCF;
                    16'hFB2D: data_out = 8'hCE;
                    16'hFB2E: data_out = 8'hCD;
                    16'hFB2F: data_out = 8'hCC;
                    16'hFB30: data_out = 8'hCB;
                    16'hFB31: data_out = 8'hCA;
                    16'hFB32: data_out = 8'hC9;
                    16'hFB33: data_out = 8'hC8;
                    16'hFB34: data_out = 8'hC7;
                    16'hFB35: data_out = 8'hC6;
                    16'hFB36: data_out = 8'hC5;
                    16'hFB37: data_out = 8'hC4;
                    16'hFB38: data_out = 8'hC3;
                    16'hFB39: data_out = 8'hC2;
                    16'hFB3A: data_out = 8'hC1;
                    16'hFB3B: data_out = 8'hC0;
                    16'hFB3C: data_out = 8'hBF;
                    16'hFB3D: data_out = 8'hBE;
                    16'hFB3E: data_out = 8'hBD;
                    16'hFB3F: data_out = 8'hBC;
                    16'hFB40: data_out = 8'hBB;
                    16'hFB41: data_out = 8'hBA;
                    16'hFB42: data_out = 8'hB9;
                    16'hFB43: data_out = 8'hB8;
                    16'hFB44: data_out = 8'hB7;
                    16'hFB45: data_out = 8'hB6;
                    16'hFB46: data_out = 8'hB5;
                    16'hFB47: data_out = 8'hB4;
                    16'hFB48: data_out = 8'hB3;
                    16'hFB49: data_out = 8'hB2;
                    16'hFB4A: data_out = 8'hB1;
                    16'hFB4B: data_out = 8'hB0;
                    16'hFB4C: data_out = 8'hAF;
                    16'hFB4D: data_out = 8'hAE;
                    16'hFB4E: data_out = 8'hAD;
                    16'hFB4F: data_out = 8'hAC;
                    16'hFB50: data_out = 8'hAB;
                    16'hFB51: data_out = 8'hAA;
                    16'hFB52: data_out = 8'hA9;
                    16'hFB53: data_out = 8'hA8;
                    16'hFB54: data_out = 8'hA7;
                    16'hFB55: data_out = 8'hA6;
                    16'hFB56: data_out = 8'hA5;
                    16'hFB57: data_out = 8'hA4;
                    16'hFB58: data_out = 8'hA3;
                    16'hFB59: data_out = 8'hA2;
                    16'hFB5A: data_out = 8'hA1;
                    16'hFB5B: data_out = 8'hA0;
                    16'hFB5C: data_out = 8'h9F;
                    16'hFB5D: data_out = 8'h9E;
                    16'hFB5E: data_out = 8'h9D;
                    16'hFB5F: data_out = 8'h9C;
                    16'hFB60: data_out = 8'h9B;
                    16'hFB61: data_out = 8'h9A;
                    16'hFB62: data_out = 8'h99;
                    16'hFB63: data_out = 8'h98;
                    16'hFB64: data_out = 8'h97;
                    16'hFB65: data_out = 8'h96;
                    16'hFB66: data_out = 8'h95;
                    16'hFB67: data_out = 8'h94;
                    16'hFB68: data_out = 8'h93;
                    16'hFB69: data_out = 8'h92;
                    16'hFB6A: data_out = 8'h91;
                    16'hFB6B: data_out = 8'h90;
                    16'hFB6C: data_out = 8'h8F;
                    16'hFB6D: data_out = 8'h8E;
                    16'hFB6E: data_out = 8'h8D;
                    16'hFB6F: data_out = 8'h8C;
                    16'hFB70: data_out = 8'h8B;
                    16'hFB71: data_out = 8'h8A;
                    16'hFB72: data_out = 8'h89;
                    16'hFB73: data_out = 8'h88;
                    16'hFB74: data_out = 8'h87;
                    16'hFB75: data_out = 8'h86;
                    16'hFB76: data_out = 8'h85;
                    16'hFB77: data_out = 8'h84;
                    16'hFB78: data_out = 8'h83;
                    16'hFB79: data_out = 8'h82;
                    16'hFB7A: data_out = 8'h81;
                    16'hFB7B: data_out = 8'h0;
                    16'hFB7C: data_out = 8'h1;
                    16'hFB7D: data_out = 8'h2;
                    16'hFB7E: data_out = 8'h3;
                    16'hFB7F: data_out = 8'h4;
                    16'hFB80: data_out = 8'hFB;
                    16'hFB81: data_out = 8'hFC;
                    16'hFB82: data_out = 8'hFD;
                    16'hFB83: data_out = 8'hFE;
                    16'hFB84: data_out = 8'hFF;
                    16'hFB85: data_out = 8'h80;
                    16'hFB86: data_out = 8'h81;
                    16'hFB87: data_out = 8'h82;
                    16'hFB88: data_out = 8'h83;
                    16'hFB89: data_out = 8'h84;
                    16'hFB8A: data_out = 8'h85;
                    16'hFB8B: data_out = 8'h86;
                    16'hFB8C: data_out = 8'h87;
                    16'hFB8D: data_out = 8'h88;
                    16'hFB8E: data_out = 8'h89;
                    16'hFB8F: data_out = 8'h8A;
                    16'hFB90: data_out = 8'h8B;
                    16'hFB91: data_out = 8'h8C;
                    16'hFB92: data_out = 8'h8D;
                    16'hFB93: data_out = 8'h8E;
                    16'hFB94: data_out = 8'h8F;
                    16'hFB95: data_out = 8'h90;
                    16'hFB96: data_out = 8'h91;
                    16'hFB97: data_out = 8'h92;
                    16'hFB98: data_out = 8'h93;
                    16'hFB99: data_out = 8'h94;
                    16'hFB9A: data_out = 8'h95;
                    16'hFB9B: data_out = 8'h96;
                    16'hFB9C: data_out = 8'h97;
                    16'hFB9D: data_out = 8'h98;
                    16'hFB9E: data_out = 8'h99;
                    16'hFB9F: data_out = 8'h9A;
                    16'hFBA0: data_out = 8'h9B;
                    16'hFBA1: data_out = 8'h9C;
                    16'hFBA2: data_out = 8'h9D;
                    16'hFBA3: data_out = 8'h9E;
                    16'hFBA4: data_out = 8'h9F;
                    16'hFBA5: data_out = 8'hA0;
                    16'hFBA6: data_out = 8'hA1;
                    16'hFBA7: data_out = 8'hA2;
                    16'hFBA8: data_out = 8'hA3;
                    16'hFBA9: data_out = 8'hA4;
                    16'hFBAA: data_out = 8'hA5;
                    16'hFBAB: data_out = 8'hA6;
                    16'hFBAC: data_out = 8'hA7;
                    16'hFBAD: data_out = 8'hA8;
                    16'hFBAE: data_out = 8'hA9;
                    16'hFBAF: data_out = 8'hAA;
                    16'hFBB0: data_out = 8'hAB;
                    16'hFBB1: data_out = 8'hAC;
                    16'hFBB2: data_out = 8'hAD;
                    16'hFBB3: data_out = 8'hAE;
                    16'hFBB4: data_out = 8'hAF;
                    16'hFBB5: data_out = 8'hB0;
                    16'hFBB6: data_out = 8'hB1;
                    16'hFBB7: data_out = 8'hB2;
                    16'hFBB8: data_out = 8'hB3;
                    16'hFBB9: data_out = 8'hB4;
                    16'hFBBA: data_out = 8'hB5;
                    16'hFBBB: data_out = 8'hB6;
                    16'hFBBC: data_out = 8'hB7;
                    16'hFBBD: data_out = 8'hB8;
                    16'hFBBE: data_out = 8'hB9;
                    16'hFBBF: data_out = 8'hBA;
                    16'hFBC0: data_out = 8'hBB;
                    16'hFBC1: data_out = 8'hBC;
                    16'hFBC2: data_out = 8'hBD;
                    16'hFBC3: data_out = 8'hBE;
                    16'hFBC4: data_out = 8'hBF;
                    16'hFBC5: data_out = 8'hC0;
                    16'hFBC6: data_out = 8'hC1;
                    16'hFBC7: data_out = 8'hC2;
                    16'hFBC8: data_out = 8'hC3;
                    16'hFBC9: data_out = 8'hC4;
                    16'hFBCA: data_out = 8'hC5;
                    16'hFBCB: data_out = 8'hC6;
                    16'hFBCC: data_out = 8'hC7;
                    16'hFBCD: data_out = 8'hC8;
                    16'hFBCE: data_out = 8'hC9;
                    16'hFBCF: data_out = 8'hCA;
                    16'hFBD0: data_out = 8'hCB;
                    16'hFBD1: data_out = 8'hCC;
                    16'hFBD2: data_out = 8'hCD;
                    16'hFBD3: data_out = 8'hCE;
                    16'hFBD4: data_out = 8'hCF;
                    16'hFBD5: data_out = 8'hD0;
                    16'hFBD6: data_out = 8'hD1;
                    16'hFBD7: data_out = 8'hD2;
                    16'hFBD8: data_out = 8'hD3;
                    16'hFBD9: data_out = 8'hD4;
                    16'hFBDA: data_out = 8'hD5;
                    16'hFBDB: data_out = 8'hD6;
                    16'hFBDC: data_out = 8'hD7;
                    16'hFBDD: data_out = 8'hD8;
                    16'hFBDE: data_out = 8'hD9;
                    16'hFBDF: data_out = 8'hDA;
                    16'hFBE0: data_out = 8'hDB;
                    16'hFBE1: data_out = 8'hDC;
                    16'hFBE2: data_out = 8'hDD;
                    16'hFBE3: data_out = 8'hDE;
                    16'hFBE4: data_out = 8'hDF;
                    16'hFBE5: data_out = 8'hE0;
                    16'hFBE6: data_out = 8'hE1;
                    16'hFBE7: data_out = 8'hE2;
                    16'hFBE8: data_out = 8'hE3;
                    16'hFBE9: data_out = 8'hE4;
                    16'hFBEA: data_out = 8'hE5;
                    16'hFBEB: data_out = 8'hE6;
                    16'hFBEC: data_out = 8'hE7;
                    16'hFBED: data_out = 8'hE8;
                    16'hFBEE: data_out = 8'hE9;
                    16'hFBEF: data_out = 8'hEA;
                    16'hFBF0: data_out = 8'hEB;
                    16'hFBF1: data_out = 8'hEC;
                    16'hFBF2: data_out = 8'hED;
                    16'hFBF3: data_out = 8'hEE;
                    16'hFBF4: data_out = 8'hEF;
                    16'hFBF5: data_out = 8'hF0;
                    16'hFBF6: data_out = 8'hF1;
                    16'hFBF7: data_out = 8'hF2;
                    16'hFBF8: data_out = 8'hF3;
                    16'hFBF9: data_out = 8'hF4;
                    16'hFBFA: data_out = 8'hF5;
                    16'hFBFB: data_out = 8'hF6;
                    16'hFBFC: data_out = 8'hF7;
                    16'hFBFD: data_out = 8'hF8;
                    16'hFBFE: data_out = 8'hF9;
                    16'hFBFF: data_out = 8'hFA;
                    16'hFC00: data_out = 8'hFC;
                    16'hFC01: data_out = 8'hFB;
                    16'hFC02: data_out = 8'hFA;
                    16'hFC03: data_out = 8'hF9;
                    16'hFC04: data_out = 8'hF8;
                    16'hFC05: data_out = 8'hF7;
                    16'hFC06: data_out = 8'hF6;
                    16'hFC07: data_out = 8'hF5;
                    16'hFC08: data_out = 8'hF4;
                    16'hFC09: data_out = 8'hF3;
                    16'hFC0A: data_out = 8'hF2;
                    16'hFC0B: data_out = 8'hF1;
                    16'hFC0C: data_out = 8'hF0;
                    16'hFC0D: data_out = 8'hEF;
                    16'hFC0E: data_out = 8'hEE;
                    16'hFC0F: data_out = 8'hED;
                    16'hFC10: data_out = 8'hEC;
                    16'hFC11: data_out = 8'hEB;
                    16'hFC12: data_out = 8'hEA;
                    16'hFC13: data_out = 8'hE9;
                    16'hFC14: data_out = 8'hE8;
                    16'hFC15: data_out = 8'hE7;
                    16'hFC16: data_out = 8'hE6;
                    16'hFC17: data_out = 8'hE5;
                    16'hFC18: data_out = 8'hE4;
                    16'hFC19: data_out = 8'hE3;
                    16'hFC1A: data_out = 8'hE2;
                    16'hFC1B: data_out = 8'hE1;
                    16'hFC1C: data_out = 8'hE0;
                    16'hFC1D: data_out = 8'hDF;
                    16'hFC1E: data_out = 8'hDE;
                    16'hFC1F: data_out = 8'hDD;
                    16'hFC20: data_out = 8'hDC;
                    16'hFC21: data_out = 8'hDB;
                    16'hFC22: data_out = 8'hDA;
                    16'hFC23: data_out = 8'hD9;
                    16'hFC24: data_out = 8'hD8;
                    16'hFC25: data_out = 8'hD7;
                    16'hFC26: data_out = 8'hD6;
                    16'hFC27: data_out = 8'hD5;
                    16'hFC28: data_out = 8'hD4;
                    16'hFC29: data_out = 8'hD3;
                    16'hFC2A: data_out = 8'hD2;
                    16'hFC2B: data_out = 8'hD1;
                    16'hFC2C: data_out = 8'hD0;
                    16'hFC2D: data_out = 8'hCF;
                    16'hFC2E: data_out = 8'hCE;
                    16'hFC2F: data_out = 8'hCD;
                    16'hFC30: data_out = 8'hCC;
                    16'hFC31: data_out = 8'hCB;
                    16'hFC32: data_out = 8'hCA;
                    16'hFC33: data_out = 8'hC9;
                    16'hFC34: data_out = 8'hC8;
                    16'hFC35: data_out = 8'hC7;
                    16'hFC36: data_out = 8'hC6;
                    16'hFC37: data_out = 8'hC5;
                    16'hFC38: data_out = 8'hC4;
                    16'hFC39: data_out = 8'hC3;
                    16'hFC3A: data_out = 8'hC2;
                    16'hFC3B: data_out = 8'hC1;
                    16'hFC3C: data_out = 8'hC0;
                    16'hFC3D: data_out = 8'hBF;
                    16'hFC3E: data_out = 8'hBE;
                    16'hFC3F: data_out = 8'hBD;
                    16'hFC40: data_out = 8'hBC;
                    16'hFC41: data_out = 8'hBB;
                    16'hFC42: data_out = 8'hBA;
                    16'hFC43: data_out = 8'hB9;
                    16'hFC44: data_out = 8'hB8;
                    16'hFC45: data_out = 8'hB7;
                    16'hFC46: data_out = 8'hB6;
                    16'hFC47: data_out = 8'hB5;
                    16'hFC48: data_out = 8'hB4;
                    16'hFC49: data_out = 8'hB3;
                    16'hFC4A: data_out = 8'hB2;
                    16'hFC4B: data_out = 8'hB1;
                    16'hFC4C: data_out = 8'hB0;
                    16'hFC4D: data_out = 8'hAF;
                    16'hFC4E: data_out = 8'hAE;
                    16'hFC4F: data_out = 8'hAD;
                    16'hFC50: data_out = 8'hAC;
                    16'hFC51: data_out = 8'hAB;
                    16'hFC52: data_out = 8'hAA;
                    16'hFC53: data_out = 8'hA9;
                    16'hFC54: data_out = 8'hA8;
                    16'hFC55: data_out = 8'hA7;
                    16'hFC56: data_out = 8'hA6;
                    16'hFC57: data_out = 8'hA5;
                    16'hFC58: data_out = 8'hA4;
                    16'hFC59: data_out = 8'hA3;
                    16'hFC5A: data_out = 8'hA2;
                    16'hFC5B: data_out = 8'hA1;
                    16'hFC5C: data_out = 8'hA0;
                    16'hFC5D: data_out = 8'h9F;
                    16'hFC5E: data_out = 8'h9E;
                    16'hFC5F: data_out = 8'h9D;
                    16'hFC60: data_out = 8'h9C;
                    16'hFC61: data_out = 8'h9B;
                    16'hFC62: data_out = 8'h9A;
                    16'hFC63: data_out = 8'h99;
                    16'hFC64: data_out = 8'h98;
                    16'hFC65: data_out = 8'h97;
                    16'hFC66: data_out = 8'h96;
                    16'hFC67: data_out = 8'h95;
                    16'hFC68: data_out = 8'h94;
                    16'hFC69: data_out = 8'h93;
                    16'hFC6A: data_out = 8'h92;
                    16'hFC6B: data_out = 8'h91;
                    16'hFC6C: data_out = 8'h90;
                    16'hFC6D: data_out = 8'h8F;
                    16'hFC6E: data_out = 8'h8E;
                    16'hFC6F: data_out = 8'h8D;
                    16'hFC70: data_out = 8'h8C;
                    16'hFC71: data_out = 8'h8B;
                    16'hFC72: data_out = 8'h8A;
                    16'hFC73: data_out = 8'h89;
                    16'hFC74: data_out = 8'h88;
                    16'hFC75: data_out = 8'h87;
                    16'hFC76: data_out = 8'h86;
                    16'hFC77: data_out = 8'h85;
                    16'hFC78: data_out = 8'h84;
                    16'hFC79: data_out = 8'h83;
                    16'hFC7A: data_out = 8'h82;
                    16'hFC7B: data_out = 8'h81;
                    16'hFC7C: data_out = 8'h0;
                    16'hFC7D: data_out = 8'h1;
                    16'hFC7E: data_out = 8'h2;
                    16'hFC7F: data_out = 8'h3;
                    16'hFC80: data_out = 8'hFC;
                    16'hFC81: data_out = 8'hFD;
                    16'hFC82: data_out = 8'hFE;
                    16'hFC83: data_out = 8'hFF;
                    16'hFC84: data_out = 8'h80;
                    16'hFC85: data_out = 8'h81;
                    16'hFC86: data_out = 8'h82;
                    16'hFC87: data_out = 8'h83;
                    16'hFC88: data_out = 8'h84;
                    16'hFC89: data_out = 8'h85;
                    16'hFC8A: data_out = 8'h86;
                    16'hFC8B: data_out = 8'h87;
                    16'hFC8C: data_out = 8'h88;
                    16'hFC8D: data_out = 8'h89;
                    16'hFC8E: data_out = 8'h8A;
                    16'hFC8F: data_out = 8'h8B;
                    16'hFC90: data_out = 8'h8C;
                    16'hFC91: data_out = 8'h8D;
                    16'hFC92: data_out = 8'h8E;
                    16'hFC93: data_out = 8'h8F;
                    16'hFC94: data_out = 8'h90;
                    16'hFC95: data_out = 8'h91;
                    16'hFC96: data_out = 8'h92;
                    16'hFC97: data_out = 8'h93;
                    16'hFC98: data_out = 8'h94;
                    16'hFC99: data_out = 8'h95;
                    16'hFC9A: data_out = 8'h96;
                    16'hFC9B: data_out = 8'h97;
                    16'hFC9C: data_out = 8'h98;
                    16'hFC9D: data_out = 8'h99;
                    16'hFC9E: data_out = 8'h9A;
                    16'hFC9F: data_out = 8'h9B;
                    16'hFCA0: data_out = 8'h9C;
                    16'hFCA1: data_out = 8'h9D;
                    16'hFCA2: data_out = 8'h9E;
                    16'hFCA3: data_out = 8'h9F;
                    16'hFCA4: data_out = 8'hA0;
                    16'hFCA5: data_out = 8'hA1;
                    16'hFCA6: data_out = 8'hA2;
                    16'hFCA7: data_out = 8'hA3;
                    16'hFCA8: data_out = 8'hA4;
                    16'hFCA9: data_out = 8'hA5;
                    16'hFCAA: data_out = 8'hA6;
                    16'hFCAB: data_out = 8'hA7;
                    16'hFCAC: data_out = 8'hA8;
                    16'hFCAD: data_out = 8'hA9;
                    16'hFCAE: data_out = 8'hAA;
                    16'hFCAF: data_out = 8'hAB;
                    16'hFCB0: data_out = 8'hAC;
                    16'hFCB1: data_out = 8'hAD;
                    16'hFCB2: data_out = 8'hAE;
                    16'hFCB3: data_out = 8'hAF;
                    16'hFCB4: data_out = 8'hB0;
                    16'hFCB5: data_out = 8'hB1;
                    16'hFCB6: data_out = 8'hB2;
                    16'hFCB7: data_out = 8'hB3;
                    16'hFCB8: data_out = 8'hB4;
                    16'hFCB9: data_out = 8'hB5;
                    16'hFCBA: data_out = 8'hB6;
                    16'hFCBB: data_out = 8'hB7;
                    16'hFCBC: data_out = 8'hB8;
                    16'hFCBD: data_out = 8'hB9;
                    16'hFCBE: data_out = 8'hBA;
                    16'hFCBF: data_out = 8'hBB;
                    16'hFCC0: data_out = 8'hBC;
                    16'hFCC1: data_out = 8'hBD;
                    16'hFCC2: data_out = 8'hBE;
                    16'hFCC3: data_out = 8'hBF;
                    16'hFCC4: data_out = 8'hC0;
                    16'hFCC5: data_out = 8'hC1;
                    16'hFCC6: data_out = 8'hC2;
                    16'hFCC7: data_out = 8'hC3;
                    16'hFCC8: data_out = 8'hC4;
                    16'hFCC9: data_out = 8'hC5;
                    16'hFCCA: data_out = 8'hC6;
                    16'hFCCB: data_out = 8'hC7;
                    16'hFCCC: data_out = 8'hC8;
                    16'hFCCD: data_out = 8'hC9;
                    16'hFCCE: data_out = 8'hCA;
                    16'hFCCF: data_out = 8'hCB;
                    16'hFCD0: data_out = 8'hCC;
                    16'hFCD1: data_out = 8'hCD;
                    16'hFCD2: data_out = 8'hCE;
                    16'hFCD3: data_out = 8'hCF;
                    16'hFCD4: data_out = 8'hD0;
                    16'hFCD5: data_out = 8'hD1;
                    16'hFCD6: data_out = 8'hD2;
                    16'hFCD7: data_out = 8'hD3;
                    16'hFCD8: data_out = 8'hD4;
                    16'hFCD9: data_out = 8'hD5;
                    16'hFCDA: data_out = 8'hD6;
                    16'hFCDB: data_out = 8'hD7;
                    16'hFCDC: data_out = 8'hD8;
                    16'hFCDD: data_out = 8'hD9;
                    16'hFCDE: data_out = 8'hDA;
                    16'hFCDF: data_out = 8'hDB;
                    16'hFCE0: data_out = 8'hDC;
                    16'hFCE1: data_out = 8'hDD;
                    16'hFCE2: data_out = 8'hDE;
                    16'hFCE3: data_out = 8'hDF;
                    16'hFCE4: data_out = 8'hE0;
                    16'hFCE5: data_out = 8'hE1;
                    16'hFCE6: data_out = 8'hE2;
                    16'hFCE7: data_out = 8'hE3;
                    16'hFCE8: data_out = 8'hE4;
                    16'hFCE9: data_out = 8'hE5;
                    16'hFCEA: data_out = 8'hE6;
                    16'hFCEB: data_out = 8'hE7;
                    16'hFCEC: data_out = 8'hE8;
                    16'hFCED: data_out = 8'hE9;
                    16'hFCEE: data_out = 8'hEA;
                    16'hFCEF: data_out = 8'hEB;
                    16'hFCF0: data_out = 8'hEC;
                    16'hFCF1: data_out = 8'hED;
                    16'hFCF2: data_out = 8'hEE;
                    16'hFCF3: data_out = 8'hEF;
                    16'hFCF4: data_out = 8'hF0;
                    16'hFCF5: data_out = 8'hF1;
                    16'hFCF6: data_out = 8'hF2;
                    16'hFCF7: data_out = 8'hF3;
                    16'hFCF8: data_out = 8'hF4;
                    16'hFCF9: data_out = 8'hF5;
                    16'hFCFA: data_out = 8'hF6;
                    16'hFCFB: data_out = 8'hF7;
                    16'hFCFC: data_out = 8'hF8;
                    16'hFCFD: data_out = 8'hF9;
                    16'hFCFE: data_out = 8'hFA;
                    16'hFCFF: data_out = 8'hFB;
                    16'hFD00: data_out = 8'hFD;
                    16'hFD01: data_out = 8'hFC;
                    16'hFD02: data_out = 8'hFB;
                    16'hFD03: data_out = 8'hFA;
                    16'hFD04: data_out = 8'hF9;
                    16'hFD05: data_out = 8'hF8;
                    16'hFD06: data_out = 8'hF7;
                    16'hFD07: data_out = 8'hF6;
                    16'hFD08: data_out = 8'hF5;
                    16'hFD09: data_out = 8'hF4;
                    16'hFD0A: data_out = 8'hF3;
                    16'hFD0B: data_out = 8'hF2;
                    16'hFD0C: data_out = 8'hF1;
                    16'hFD0D: data_out = 8'hF0;
                    16'hFD0E: data_out = 8'hEF;
                    16'hFD0F: data_out = 8'hEE;
                    16'hFD10: data_out = 8'hED;
                    16'hFD11: data_out = 8'hEC;
                    16'hFD12: data_out = 8'hEB;
                    16'hFD13: data_out = 8'hEA;
                    16'hFD14: data_out = 8'hE9;
                    16'hFD15: data_out = 8'hE8;
                    16'hFD16: data_out = 8'hE7;
                    16'hFD17: data_out = 8'hE6;
                    16'hFD18: data_out = 8'hE5;
                    16'hFD19: data_out = 8'hE4;
                    16'hFD1A: data_out = 8'hE3;
                    16'hFD1B: data_out = 8'hE2;
                    16'hFD1C: data_out = 8'hE1;
                    16'hFD1D: data_out = 8'hE0;
                    16'hFD1E: data_out = 8'hDF;
                    16'hFD1F: data_out = 8'hDE;
                    16'hFD20: data_out = 8'hDD;
                    16'hFD21: data_out = 8'hDC;
                    16'hFD22: data_out = 8'hDB;
                    16'hFD23: data_out = 8'hDA;
                    16'hFD24: data_out = 8'hD9;
                    16'hFD25: data_out = 8'hD8;
                    16'hFD26: data_out = 8'hD7;
                    16'hFD27: data_out = 8'hD6;
                    16'hFD28: data_out = 8'hD5;
                    16'hFD29: data_out = 8'hD4;
                    16'hFD2A: data_out = 8'hD3;
                    16'hFD2B: data_out = 8'hD2;
                    16'hFD2C: data_out = 8'hD1;
                    16'hFD2D: data_out = 8'hD0;
                    16'hFD2E: data_out = 8'hCF;
                    16'hFD2F: data_out = 8'hCE;
                    16'hFD30: data_out = 8'hCD;
                    16'hFD31: data_out = 8'hCC;
                    16'hFD32: data_out = 8'hCB;
                    16'hFD33: data_out = 8'hCA;
                    16'hFD34: data_out = 8'hC9;
                    16'hFD35: data_out = 8'hC8;
                    16'hFD36: data_out = 8'hC7;
                    16'hFD37: data_out = 8'hC6;
                    16'hFD38: data_out = 8'hC5;
                    16'hFD39: data_out = 8'hC4;
                    16'hFD3A: data_out = 8'hC3;
                    16'hFD3B: data_out = 8'hC2;
                    16'hFD3C: data_out = 8'hC1;
                    16'hFD3D: data_out = 8'hC0;
                    16'hFD3E: data_out = 8'hBF;
                    16'hFD3F: data_out = 8'hBE;
                    16'hFD40: data_out = 8'hBD;
                    16'hFD41: data_out = 8'hBC;
                    16'hFD42: data_out = 8'hBB;
                    16'hFD43: data_out = 8'hBA;
                    16'hFD44: data_out = 8'hB9;
                    16'hFD45: data_out = 8'hB8;
                    16'hFD46: data_out = 8'hB7;
                    16'hFD47: data_out = 8'hB6;
                    16'hFD48: data_out = 8'hB5;
                    16'hFD49: data_out = 8'hB4;
                    16'hFD4A: data_out = 8'hB3;
                    16'hFD4B: data_out = 8'hB2;
                    16'hFD4C: data_out = 8'hB1;
                    16'hFD4D: data_out = 8'hB0;
                    16'hFD4E: data_out = 8'hAF;
                    16'hFD4F: data_out = 8'hAE;
                    16'hFD50: data_out = 8'hAD;
                    16'hFD51: data_out = 8'hAC;
                    16'hFD52: data_out = 8'hAB;
                    16'hFD53: data_out = 8'hAA;
                    16'hFD54: data_out = 8'hA9;
                    16'hFD55: data_out = 8'hA8;
                    16'hFD56: data_out = 8'hA7;
                    16'hFD57: data_out = 8'hA6;
                    16'hFD58: data_out = 8'hA5;
                    16'hFD59: data_out = 8'hA4;
                    16'hFD5A: data_out = 8'hA3;
                    16'hFD5B: data_out = 8'hA2;
                    16'hFD5C: data_out = 8'hA1;
                    16'hFD5D: data_out = 8'hA0;
                    16'hFD5E: data_out = 8'h9F;
                    16'hFD5F: data_out = 8'h9E;
                    16'hFD60: data_out = 8'h9D;
                    16'hFD61: data_out = 8'h9C;
                    16'hFD62: data_out = 8'h9B;
                    16'hFD63: data_out = 8'h9A;
                    16'hFD64: data_out = 8'h99;
                    16'hFD65: data_out = 8'h98;
                    16'hFD66: data_out = 8'h97;
                    16'hFD67: data_out = 8'h96;
                    16'hFD68: data_out = 8'h95;
                    16'hFD69: data_out = 8'h94;
                    16'hFD6A: data_out = 8'h93;
                    16'hFD6B: data_out = 8'h92;
                    16'hFD6C: data_out = 8'h91;
                    16'hFD6D: data_out = 8'h90;
                    16'hFD6E: data_out = 8'h8F;
                    16'hFD6F: data_out = 8'h8E;
                    16'hFD70: data_out = 8'h8D;
                    16'hFD71: data_out = 8'h8C;
                    16'hFD72: data_out = 8'h8B;
                    16'hFD73: data_out = 8'h8A;
                    16'hFD74: data_out = 8'h89;
                    16'hFD75: data_out = 8'h88;
                    16'hFD76: data_out = 8'h87;
                    16'hFD77: data_out = 8'h86;
                    16'hFD78: data_out = 8'h85;
                    16'hFD79: data_out = 8'h84;
                    16'hFD7A: data_out = 8'h83;
                    16'hFD7B: data_out = 8'h82;
                    16'hFD7C: data_out = 8'h81;
                    16'hFD7D: data_out = 8'h0;
                    16'hFD7E: data_out = 8'h1;
                    16'hFD7F: data_out = 8'h2;
                    16'hFD80: data_out = 8'hFD;
                    16'hFD81: data_out = 8'hFE;
                    16'hFD82: data_out = 8'hFF;
                    16'hFD83: data_out = 8'h80;
                    16'hFD84: data_out = 8'h81;
                    16'hFD85: data_out = 8'h82;
                    16'hFD86: data_out = 8'h83;
                    16'hFD87: data_out = 8'h84;
                    16'hFD88: data_out = 8'h85;
                    16'hFD89: data_out = 8'h86;
                    16'hFD8A: data_out = 8'h87;
                    16'hFD8B: data_out = 8'h88;
                    16'hFD8C: data_out = 8'h89;
                    16'hFD8D: data_out = 8'h8A;
                    16'hFD8E: data_out = 8'h8B;
                    16'hFD8F: data_out = 8'h8C;
                    16'hFD90: data_out = 8'h8D;
                    16'hFD91: data_out = 8'h8E;
                    16'hFD92: data_out = 8'h8F;
                    16'hFD93: data_out = 8'h90;
                    16'hFD94: data_out = 8'h91;
                    16'hFD95: data_out = 8'h92;
                    16'hFD96: data_out = 8'h93;
                    16'hFD97: data_out = 8'h94;
                    16'hFD98: data_out = 8'h95;
                    16'hFD99: data_out = 8'h96;
                    16'hFD9A: data_out = 8'h97;
                    16'hFD9B: data_out = 8'h98;
                    16'hFD9C: data_out = 8'h99;
                    16'hFD9D: data_out = 8'h9A;
                    16'hFD9E: data_out = 8'h9B;
                    16'hFD9F: data_out = 8'h9C;
                    16'hFDA0: data_out = 8'h9D;
                    16'hFDA1: data_out = 8'h9E;
                    16'hFDA2: data_out = 8'h9F;
                    16'hFDA3: data_out = 8'hA0;
                    16'hFDA4: data_out = 8'hA1;
                    16'hFDA5: data_out = 8'hA2;
                    16'hFDA6: data_out = 8'hA3;
                    16'hFDA7: data_out = 8'hA4;
                    16'hFDA8: data_out = 8'hA5;
                    16'hFDA9: data_out = 8'hA6;
                    16'hFDAA: data_out = 8'hA7;
                    16'hFDAB: data_out = 8'hA8;
                    16'hFDAC: data_out = 8'hA9;
                    16'hFDAD: data_out = 8'hAA;
                    16'hFDAE: data_out = 8'hAB;
                    16'hFDAF: data_out = 8'hAC;
                    16'hFDB0: data_out = 8'hAD;
                    16'hFDB1: data_out = 8'hAE;
                    16'hFDB2: data_out = 8'hAF;
                    16'hFDB3: data_out = 8'hB0;
                    16'hFDB4: data_out = 8'hB1;
                    16'hFDB5: data_out = 8'hB2;
                    16'hFDB6: data_out = 8'hB3;
                    16'hFDB7: data_out = 8'hB4;
                    16'hFDB8: data_out = 8'hB5;
                    16'hFDB9: data_out = 8'hB6;
                    16'hFDBA: data_out = 8'hB7;
                    16'hFDBB: data_out = 8'hB8;
                    16'hFDBC: data_out = 8'hB9;
                    16'hFDBD: data_out = 8'hBA;
                    16'hFDBE: data_out = 8'hBB;
                    16'hFDBF: data_out = 8'hBC;
                    16'hFDC0: data_out = 8'hBD;
                    16'hFDC1: data_out = 8'hBE;
                    16'hFDC2: data_out = 8'hBF;
                    16'hFDC3: data_out = 8'hC0;
                    16'hFDC4: data_out = 8'hC1;
                    16'hFDC5: data_out = 8'hC2;
                    16'hFDC6: data_out = 8'hC3;
                    16'hFDC7: data_out = 8'hC4;
                    16'hFDC8: data_out = 8'hC5;
                    16'hFDC9: data_out = 8'hC6;
                    16'hFDCA: data_out = 8'hC7;
                    16'hFDCB: data_out = 8'hC8;
                    16'hFDCC: data_out = 8'hC9;
                    16'hFDCD: data_out = 8'hCA;
                    16'hFDCE: data_out = 8'hCB;
                    16'hFDCF: data_out = 8'hCC;
                    16'hFDD0: data_out = 8'hCD;
                    16'hFDD1: data_out = 8'hCE;
                    16'hFDD2: data_out = 8'hCF;
                    16'hFDD3: data_out = 8'hD0;
                    16'hFDD4: data_out = 8'hD1;
                    16'hFDD5: data_out = 8'hD2;
                    16'hFDD6: data_out = 8'hD3;
                    16'hFDD7: data_out = 8'hD4;
                    16'hFDD8: data_out = 8'hD5;
                    16'hFDD9: data_out = 8'hD6;
                    16'hFDDA: data_out = 8'hD7;
                    16'hFDDB: data_out = 8'hD8;
                    16'hFDDC: data_out = 8'hD9;
                    16'hFDDD: data_out = 8'hDA;
                    16'hFDDE: data_out = 8'hDB;
                    16'hFDDF: data_out = 8'hDC;
                    16'hFDE0: data_out = 8'hDD;
                    16'hFDE1: data_out = 8'hDE;
                    16'hFDE2: data_out = 8'hDF;
                    16'hFDE3: data_out = 8'hE0;
                    16'hFDE4: data_out = 8'hE1;
                    16'hFDE5: data_out = 8'hE2;
                    16'hFDE6: data_out = 8'hE3;
                    16'hFDE7: data_out = 8'hE4;
                    16'hFDE8: data_out = 8'hE5;
                    16'hFDE9: data_out = 8'hE6;
                    16'hFDEA: data_out = 8'hE7;
                    16'hFDEB: data_out = 8'hE8;
                    16'hFDEC: data_out = 8'hE9;
                    16'hFDED: data_out = 8'hEA;
                    16'hFDEE: data_out = 8'hEB;
                    16'hFDEF: data_out = 8'hEC;
                    16'hFDF0: data_out = 8'hED;
                    16'hFDF1: data_out = 8'hEE;
                    16'hFDF2: data_out = 8'hEF;
                    16'hFDF3: data_out = 8'hF0;
                    16'hFDF4: data_out = 8'hF1;
                    16'hFDF5: data_out = 8'hF2;
                    16'hFDF6: data_out = 8'hF3;
                    16'hFDF7: data_out = 8'hF4;
                    16'hFDF8: data_out = 8'hF5;
                    16'hFDF9: data_out = 8'hF6;
                    16'hFDFA: data_out = 8'hF7;
                    16'hFDFB: data_out = 8'hF8;
                    16'hFDFC: data_out = 8'hF9;
                    16'hFDFD: data_out = 8'hFA;
                    16'hFDFE: data_out = 8'hFB;
                    16'hFDFF: data_out = 8'hFC;
                    16'hFE00: data_out = 8'hFE;
                    16'hFE01: data_out = 8'hFD;
                    16'hFE02: data_out = 8'hFC;
                    16'hFE03: data_out = 8'hFB;
                    16'hFE04: data_out = 8'hFA;
                    16'hFE05: data_out = 8'hF9;
                    16'hFE06: data_out = 8'hF8;
                    16'hFE07: data_out = 8'hF7;
                    16'hFE08: data_out = 8'hF6;
                    16'hFE09: data_out = 8'hF5;
                    16'hFE0A: data_out = 8'hF4;
                    16'hFE0B: data_out = 8'hF3;
                    16'hFE0C: data_out = 8'hF2;
                    16'hFE0D: data_out = 8'hF1;
                    16'hFE0E: data_out = 8'hF0;
                    16'hFE0F: data_out = 8'hEF;
                    16'hFE10: data_out = 8'hEE;
                    16'hFE11: data_out = 8'hED;
                    16'hFE12: data_out = 8'hEC;
                    16'hFE13: data_out = 8'hEB;
                    16'hFE14: data_out = 8'hEA;
                    16'hFE15: data_out = 8'hE9;
                    16'hFE16: data_out = 8'hE8;
                    16'hFE17: data_out = 8'hE7;
                    16'hFE18: data_out = 8'hE6;
                    16'hFE19: data_out = 8'hE5;
                    16'hFE1A: data_out = 8'hE4;
                    16'hFE1B: data_out = 8'hE3;
                    16'hFE1C: data_out = 8'hE2;
                    16'hFE1D: data_out = 8'hE1;
                    16'hFE1E: data_out = 8'hE0;
                    16'hFE1F: data_out = 8'hDF;
                    16'hFE20: data_out = 8'hDE;
                    16'hFE21: data_out = 8'hDD;
                    16'hFE22: data_out = 8'hDC;
                    16'hFE23: data_out = 8'hDB;
                    16'hFE24: data_out = 8'hDA;
                    16'hFE25: data_out = 8'hD9;
                    16'hFE26: data_out = 8'hD8;
                    16'hFE27: data_out = 8'hD7;
                    16'hFE28: data_out = 8'hD6;
                    16'hFE29: data_out = 8'hD5;
                    16'hFE2A: data_out = 8'hD4;
                    16'hFE2B: data_out = 8'hD3;
                    16'hFE2C: data_out = 8'hD2;
                    16'hFE2D: data_out = 8'hD1;
                    16'hFE2E: data_out = 8'hD0;
                    16'hFE2F: data_out = 8'hCF;
                    16'hFE30: data_out = 8'hCE;
                    16'hFE31: data_out = 8'hCD;
                    16'hFE32: data_out = 8'hCC;
                    16'hFE33: data_out = 8'hCB;
                    16'hFE34: data_out = 8'hCA;
                    16'hFE35: data_out = 8'hC9;
                    16'hFE36: data_out = 8'hC8;
                    16'hFE37: data_out = 8'hC7;
                    16'hFE38: data_out = 8'hC6;
                    16'hFE39: data_out = 8'hC5;
                    16'hFE3A: data_out = 8'hC4;
                    16'hFE3B: data_out = 8'hC3;
                    16'hFE3C: data_out = 8'hC2;
                    16'hFE3D: data_out = 8'hC1;
                    16'hFE3E: data_out = 8'hC0;
                    16'hFE3F: data_out = 8'hBF;
                    16'hFE40: data_out = 8'hBE;
                    16'hFE41: data_out = 8'hBD;
                    16'hFE42: data_out = 8'hBC;
                    16'hFE43: data_out = 8'hBB;
                    16'hFE44: data_out = 8'hBA;
                    16'hFE45: data_out = 8'hB9;
                    16'hFE46: data_out = 8'hB8;
                    16'hFE47: data_out = 8'hB7;
                    16'hFE48: data_out = 8'hB6;
                    16'hFE49: data_out = 8'hB5;
                    16'hFE4A: data_out = 8'hB4;
                    16'hFE4B: data_out = 8'hB3;
                    16'hFE4C: data_out = 8'hB2;
                    16'hFE4D: data_out = 8'hB1;
                    16'hFE4E: data_out = 8'hB0;
                    16'hFE4F: data_out = 8'hAF;
                    16'hFE50: data_out = 8'hAE;
                    16'hFE51: data_out = 8'hAD;
                    16'hFE52: data_out = 8'hAC;
                    16'hFE53: data_out = 8'hAB;
                    16'hFE54: data_out = 8'hAA;
                    16'hFE55: data_out = 8'hA9;
                    16'hFE56: data_out = 8'hA8;
                    16'hFE57: data_out = 8'hA7;
                    16'hFE58: data_out = 8'hA6;
                    16'hFE59: data_out = 8'hA5;
                    16'hFE5A: data_out = 8'hA4;
                    16'hFE5B: data_out = 8'hA3;
                    16'hFE5C: data_out = 8'hA2;
                    16'hFE5D: data_out = 8'hA1;
                    16'hFE5E: data_out = 8'hA0;
                    16'hFE5F: data_out = 8'h9F;
                    16'hFE60: data_out = 8'h9E;
                    16'hFE61: data_out = 8'h9D;
                    16'hFE62: data_out = 8'h9C;
                    16'hFE63: data_out = 8'h9B;
                    16'hFE64: data_out = 8'h9A;
                    16'hFE65: data_out = 8'h99;
                    16'hFE66: data_out = 8'h98;
                    16'hFE67: data_out = 8'h97;
                    16'hFE68: data_out = 8'h96;
                    16'hFE69: data_out = 8'h95;
                    16'hFE6A: data_out = 8'h94;
                    16'hFE6B: data_out = 8'h93;
                    16'hFE6C: data_out = 8'h92;
                    16'hFE6D: data_out = 8'h91;
                    16'hFE6E: data_out = 8'h90;
                    16'hFE6F: data_out = 8'h8F;
                    16'hFE70: data_out = 8'h8E;
                    16'hFE71: data_out = 8'h8D;
                    16'hFE72: data_out = 8'h8C;
                    16'hFE73: data_out = 8'h8B;
                    16'hFE74: data_out = 8'h8A;
                    16'hFE75: data_out = 8'h89;
                    16'hFE76: data_out = 8'h88;
                    16'hFE77: data_out = 8'h87;
                    16'hFE78: data_out = 8'h86;
                    16'hFE79: data_out = 8'h85;
                    16'hFE7A: data_out = 8'h84;
                    16'hFE7B: data_out = 8'h83;
                    16'hFE7C: data_out = 8'h82;
                    16'hFE7D: data_out = 8'h81;
                    16'hFE7E: data_out = 8'h0;
                    16'hFE7F: data_out = 8'h1;
                    16'hFE80: data_out = 8'hFE;
                    16'hFE81: data_out = 8'hFF;
                    16'hFE82: data_out = 8'h80;
                    16'hFE83: data_out = 8'h81;
                    16'hFE84: data_out = 8'h82;
                    16'hFE85: data_out = 8'h83;
                    16'hFE86: data_out = 8'h84;
                    16'hFE87: data_out = 8'h85;
                    16'hFE88: data_out = 8'h86;
                    16'hFE89: data_out = 8'h87;
                    16'hFE8A: data_out = 8'h88;
                    16'hFE8B: data_out = 8'h89;
                    16'hFE8C: data_out = 8'h8A;
                    16'hFE8D: data_out = 8'h8B;
                    16'hFE8E: data_out = 8'h8C;
                    16'hFE8F: data_out = 8'h8D;
                    16'hFE90: data_out = 8'h8E;
                    16'hFE91: data_out = 8'h8F;
                    16'hFE92: data_out = 8'h90;
                    16'hFE93: data_out = 8'h91;
                    16'hFE94: data_out = 8'h92;
                    16'hFE95: data_out = 8'h93;
                    16'hFE96: data_out = 8'h94;
                    16'hFE97: data_out = 8'h95;
                    16'hFE98: data_out = 8'h96;
                    16'hFE99: data_out = 8'h97;
                    16'hFE9A: data_out = 8'h98;
                    16'hFE9B: data_out = 8'h99;
                    16'hFE9C: data_out = 8'h9A;
                    16'hFE9D: data_out = 8'h9B;
                    16'hFE9E: data_out = 8'h9C;
                    16'hFE9F: data_out = 8'h9D;
                    16'hFEA0: data_out = 8'h9E;
                    16'hFEA1: data_out = 8'h9F;
                    16'hFEA2: data_out = 8'hA0;
                    16'hFEA3: data_out = 8'hA1;
                    16'hFEA4: data_out = 8'hA2;
                    16'hFEA5: data_out = 8'hA3;
                    16'hFEA6: data_out = 8'hA4;
                    16'hFEA7: data_out = 8'hA5;
                    16'hFEA8: data_out = 8'hA6;
                    16'hFEA9: data_out = 8'hA7;
                    16'hFEAA: data_out = 8'hA8;
                    16'hFEAB: data_out = 8'hA9;
                    16'hFEAC: data_out = 8'hAA;
                    16'hFEAD: data_out = 8'hAB;
                    16'hFEAE: data_out = 8'hAC;
                    16'hFEAF: data_out = 8'hAD;
                    16'hFEB0: data_out = 8'hAE;
                    16'hFEB1: data_out = 8'hAF;
                    16'hFEB2: data_out = 8'hB0;
                    16'hFEB3: data_out = 8'hB1;
                    16'hFEB4: data_out = 8'hB2;
                    16'hFEB5: data_out = 8'hB3;
                    16'hFEB6: data_out = 8'hB4;
                    16'hFEB7: data_out = 8'hB5;
                    16'hFEB8: data_out = 8'hB6;
                    16'hFEB9: data_out = 8'hB7;
                    16'hFEBA: data_out = 8'hB8;
                    16'hFEBB: data_out = 8'hB9;
                    16'hFEBC: data_out = 8'hBA;
                    16'hFEBD: data_out = 8'hBB;
                    16'hFEBE: data_out = 8'hBC;
                    16'hFEBF: data_out = 8'hBD;
                    16'hFEC0: data_out = 8'hBE;
                    16'hFEC1: data_out = 8'hBF;
                    16'hFEC2: data_out = 8'hC0;
                    16'hFEC3: data_out = 8'hC1;
                    16'hFEC4: data_out = 8'hC2;
                    16'hFEC5: data_out = 8'hC3;
                    16'hFEC6: data_out = 8'hC4;
                    16'hFEC7: data_out = 8'hC5;
                    16'hFEC8: data_out = 8'hC6;
                    16'hFEC9: data_out = 8'hC7;
                    16'hFECA: data_out = 8'hC8;
                    16'hFECB: data_out = 8'hC9;
                    16'hFECC: data_out = 8'hCA;
                    16'hFECD: data_out = 8'hCB;
                    16'hFECE: data_out = 8'hCC;
                    16'hFECF: data_out = 8'hCD;
                    16'hFED0: data_out = 8'hCE;
                    16'hFED1: data_out = 8'hCF;
                    16'hFED2: data_out = 8'hD0;
                    16'hFED3: data_out = 8'hD1;
                    16'hFED4: data_out = 8'hD2;
                    16'hFED5: data_out = 8'hD3;
                    16'hFED6: data_out = 8'hD4;
                    16'hFED7: data_out = 8'hD5;
                    16'hFED8: data_out = 8'hD6;
                    16'hFED9: data_out = 8'hD7;
                    16'hFEDA: data_out = 8'hD8;
                    16'hFEDB: data_out = 8'hD9;
                    16'hFEDC: data_out = 8'hDA;
                    16'hFEDD: data_out = 8'hDB;
                    16'hFEDE: data_out = 8'hDC;
                    16'hFEDF: data_out = 8'hDD;
                    16'hFEE0: data_out = 8'hDE;
                    16'hFEE1: data_out = 8'hDF;
                    16'hFEE2: data_out = 8'hE0;
                    16'hFEE3: data_out = 8'hE1;
                    16'hFEE4: data_out = 8'hE2;
                    16'hFEE5: data_out = 8'hE3;
                    16'hFEE6: data_out = 8'hE4;
                    16'hFEE7: data_out = 8'hE5;
                    16'hFEE8: data_out = 8'hE6;
                    16'hFEE9: data_out = 8'hE7;
                    16'hFEEA: data_out = 8'hE8;
                    16'hFEEB: data_out = 8'hE9;
                    16'hFEEC: data_out = 8'hEA;
                    16'hFEED: data_out = 8'hEB;
                    16'hFEEE: data_out = 8'hEC;
                    16'hFEEF: data_out = 8'hED;
                    16'hFEF0: data_out = 8'hEE;
                    16'hFEF1: data_out = 8'hEF;
                    16'hFEF2: data_out = 8'hF0;
                    16'hFEF3: data_out = 8'hF1;
                    16'hFEF4: data_out = 8'hF2;
                    16'hFEF5: data_out = 8'hF3;
                    16'hFEF6: data_out = 8'hF4;
                    16'hFEF7: data_out = 8'hF5;
                    16'hFEF8: data_out = 8'hF6;
                    16'hFEF9: data_out = 8'hF7;
                    16'hFEFA: data_out = 8'hF8;
                    16'hFEFB: data_out = 8'hF9;
                    16'hFEFC: data_out = 8'hFA;
                    16'hFEFD: data_out = 8'hFB;
                    16'hFEFE: data_out = 8'hFC;
                    16'hFEFF: data_out = 8'hFD;
                    16'hFF00: data_out = 8'hFF;
                    16'hFF01: data_out = 8'hFE;
                    16'hFF02: data_out = 8'hFD;
                    16'hFF03: data_out = 8'hFC;
                    16'hFF04: data_out = 8'hFB;
                    16'hFF05: data_out = 8'hFA;
                    16'hFF06: data_out = 8'hF9;
                    16'hFF07: data_out = 8'hF8;
                    16'hFF08: data_out = 8'hF7;
                    16'hFF09: data_out = 8'hF6;
                    16'hFF0A: data_out = 8'hF5;
                    16'hFF0B: data_out = 8'hF4;
                    16'hFF0C: data_out = 8'hF3;
                    16'hFF0D: data_out = 8'hF2;
                    16'hFF0E: data_out = 8'hF1;
                    16'hFF0F: data_out = 8'hF0;
                    16'hFF10: data_out = 8'hEF;
                    16'hFF11: data_out = 8'hEE;
                    16'hFF12: data_out = 8'hED;
                    16'hFF13: data_out = 8'hEC;
                    16'hFF14: data_out = 8'hEB;
                    16'hFF15: data_out = 8'hEA;
                    16'hFF16: data_out = 8'hE9;
                    16'hFF17: data_out = 8'hE8;
                    16'hFF18: data_out = 8'hE7;
                    16'hFF19: data_out = 8'hE6;
                    16'hFF1A: data_out = 8'hE5;
                    16'hFF1B: data_out = 8'hE4;
                    16'hFF1C: data_out = 8'hE3;
                    16'hFF1D: data_out = 8'hE2;
                    16'hFF1E: data_out = 8'hE1;
                    16'hFF1F: data_out = 8'hE0;
                    16'hFF20: data_out = 8'hDF;
                    16'hFF21: data_out = 8'hDE;
                    16'hFF22: data_out = 8'hDD;
                    16'hFF23: data_out = 8'hDC;
                    16'hFF24: data_out = 8'hDB;
                    16'hFF25: data_out = 8'hDA;
                    16'hFF26: data_out = 8'hD9;
                    16'hFF27: data_out = 8'hD8;
                    16'hFF28: data_out = 8'hD7;
                    16'hFF29: data_out = 8'hD6;
                    16'hFF2A: data_out = 8'hD5;
                    16'hFF2B: data_out = 8'hD4;
                    16'hFF2C: data_out = 8'hD3;
                    16'hFF2D: data_out = 8'hD2;
                    16'hFF2E: data_out = 8'hD1;
                    16'hFF2F: data_out = 8'hD0;
                    16'hFF30: data_out = 8'hCF;
                    16'hFF31: data_out = 8'hCE;
                    16'hFF32: data_out = 8'hCD;
                    16'hFF33: data_out = 8'hCC;
                    16'hFF34: data_out = 8'hCB;
                    16'hFF35: data_out = 8'hCA;
                    16'hFF36: data_out = 8'hC9;
                    16'hFF37: data_out = 8'hC8;
                    16'hFF38: data_out = 8'hC7;
                    16'hFF39: data_out = 8'hC6;
                    16'hFF3A: data_out = 8'hC5;
                    16'hFF3B: data_out = 8'hC4;
                    16'hFF3C: data_out = 8'hC3;
                    16'hFF3D: data_out = 8'hC2;
                    16'hFF3E: data_out = 8'hC1;
                    16'hFF3F: data_out = 8'hC0;
                    16'hFF40: data_out = 8'hBF;
                    16'hFF41: data_out = 8'hBE;
                    16'hFF42: data_out = 8'hBD;
                    16'hFF43: data_out = 8'hBC;
                    16'hFF44: data_out = 8'hBB;
                    16'hFF45: data_out = 8'hBA;
                    16'hFF46: data_out = 8'hB9;
                    16'hFF47: data_out = 8'hB8;
                    16'hFF48: data_out = 8'hB7;
                    16'hFF49: data_out = 8'hB6;
                    16'hFF4A: data_out = 8'hB5;
                    16'hFF4B: data_out = 8'hB4;
                    16'hFF4C: data_out = 8'hB3;
                    16'hFF4D: data_out = 8'hB2;
                    16'hFF4E: data_out = 8'hB1;
                    16'hFF4F: data_out = 8'hB0;
                    16'hFF50: data_out = 8'hAF;
                    16'hFF51: data_out = 8'hAE;
                    16'hFF52: data_out = 8'hAD;
                    16'hFF53: data_out = 8'hAC;
                    16'hFF54: data_out = 8'hAB;
                    16'hFF55: data_out = 8'hAA;
                    16'hFF56: data_out = 8'hA9;
                    16'hFF57: data_out = 8'hA8;
                    16'hFF58: data_out = 8'hA7;
                    16'hFF59: data_out = 8'hA6;
                    16'hFF5A: data_out = 8'hA5;
                    16'hFF5B: data_out = 8'hA4;
                    16'hFF5C: data_out = 8'hA3;
                    16'hFF5D: data_out = 8'hA2;
                    16'hFF5E: data_out = 8'hA1;
                    16'hFF5F: data_out = 8'hA0;
                    16'hFF60: data_out = 8'h9F;
                    16'hFF61: data_out = 8'h9E;
                    16'hFF62: data_out = 8'h9D;
                    16'hFF63: data_out = 8'h9C;
                    16'hFF64: data_out = 8'h9B;
                    16'hFF65: data_out = 8'h9A;
                    16'hFF66: data_out = 8'h99;
                    16'hFF67: data_out = 8'h98;
                    16'hFF68: data_out = 8'h97;
                    16'hFF69: data_out = 8'h96;
                    16'hFF6A: data_out = 8'h95;
                    16'hFF6B: data_out = 8'h94;
                    16'hFF6C: data_out = 8'h93;
                    16'hFF6D: data_out = 8'h92;
                    16'hFF6E: data_out = 8'h91;
                    16'hFF6F: data_out = 8'h90;
                    16'hFF70: data_out = 8'h8F;
                    16'hFF71: data_out = 8'h8E;
                    16'hFF72: data_out = 8'h8D;
                    16'hFF73: data_out = 8'h8C;
                    16'hFF74: data_out = 8'h8B;
                    16'hFF75: data_out = 8'h8A;
                    16'hFF76: data_out = 8'h89;
                    16'hFF77: data_out = 8'h88;
                    16'hFF78: data_out = 8'h87;
                    16'hFF79: data_out = 8'h86;
                    16'hFF7A: data_out = 8'h85;
                    16'hFF7B: data_out = 8'h84;
                    16'hFF7C: data_out = 8'h83;
                    16'hFF7D: data_out = 8'h82;
                    16'hFF7E: data_out = 8'h81;
                    16'hFF7F: data_out = 8'h0;
                    16'hFF80: data_out = 8'hFF;
                    16'hFF81: data_out = 8'h80;
                    16'hFF82: data_out = 8'h81;
                    16'hFF83: data_out = 8'h82;
                    16'hFF84: data_out = 8'h83;
                    16'hFF85: data_out = 8'h84;
                    16'hFF86: data_out = 8'h85;
                    16'hFF87: data_out = 8'h86;
                    16'hFF88: data_out = 8'h87;
                    16'hFF89: data_out = 8'h88;
                    16'hFF8A: data_out = 8'h89;
                    16'hFF8B: data_out = 8'h8A;
                    16'hFF8C: data_out = 8'h8B;
                    16'hFF8D: data_out = 8'h8C;
                    16'hFF8E: data_out = 8'h8D;
                    16'hFF8F: data_out = 8'h8E;
                    16'hFF90: data_out = 8'h8F;
                    16'hFF91: data_out = 8'h90;
                    16'hFF92: data_out = 8'h91;
                    16'hFF93: data_out = 8'h92;
                    16'hFF94: data_out = 8'h93;
                    16'hFF95: data_out = 8'h94;
                    16'hFF96: data_out = 8'h95;
                    16'hFF97: data_out = 8'h96;
                    16'hFF98: data_out = 8'h97;
                    16'hFF99: data_out = 8'h98;
                    16'hFF9A: data_out = 8'h99;
                    16'hFF9B: data_out = 8'h9A;
                    16'hFF9C: data_out = 8'h9B;
                    16'hFF9D: data_out = 8'h9C;
                    16'hFF9E: data_out = 8'h9D;
                    16'hFF9F: data_out = 8'h9E;
                    16'hFFA0: data_out = 8'h9F;
                    16'hFFA1: data_out = 8'hA0;
                    16'hFFA2: data_out = 8'hA1;
                    16'hFFA3: data_out = 8'hA2;
                    16'hFFA4: data_out = 8'hA3;
                    16'hFFA5: data_out = 8'hA4;
                    16'hFFA6: data_out = 8'hA5;
                    16'hFFA7: data_out = 8'hA6;
                    16'hFFA8: data_out = 8'hA7;
                    16'hFFA9: data_out = 8'hA8;
                    16'hFFAA: data_out = 8'hA9;
                    16'hFFAB: data_out = 8'hAA;
                    16'hFFAC: data_out = 8'hAB;
                    16'hFFAD: data_out = 8'hAC;
                    16'hFFAE: data_out = 8'hAD;
                    16'hFFAF: data_out = 8'hAE;
                    16'hFFB0: data_out = 8'hAF;
                    16'hFFB1: data_out = 8'hB0;
                    16'hFFB2: data_out = 8'hB1;
                    16'hFFB3: data_out = 8'hB2;
                    16'hFFB4: data_out = 8'hB3;
                    16'hFFB5: data_out = 8'hB4;
                    16'hFFB6: data_out = 8'hB5;
                    16'hFFB7: data_out = 8'hB6;
                    16'hFFB8: data_out = 8'hB7;
                    16'hFFB9: data_out = 8'hB8;
                    16'hFFBA: data_out = 8'hB9;
                    16'hFFBB: data_out = 8'hBA;
                    16'hFFBC: data_out = 8'hBB;
                    16'hFFBD: data_out = 8'hBC;
                    16'hFFBE: data_out = 8'hBD;
                    16'hFFBF: data_out = 8'hBE;
                    16'hFFC0: data_out = 8'hBF;
                    16'hFFC1: data_out = 8'hC0;
                    16'hFFC2: data_out = 8'hC1;
                    16'hFFC3: data_out = 8'hC2;
                    16'hFFC4: data_out = 8'hC3;
                    16'hFFC5: data_out = 8'hC4;
                    16'hFFC6: data_out = 8'hC5;
                    16'hFFC7: data_out = 8'hC6;
                    16'hFFC8: data_out = 8'hC7;
                    16'hFFC9: data_out = 8'hC8;
                    16'hFFCA: data_out = 8'hC9;
                    16'hFFCB: data_out = 8'hCA;
                    16'hFFCC: data_out = 8'hCB;
                    16'hFFCD: data_out = 8'hCC;
                    16'hFFCE: data_out = 8'hCD;
                    16'hFFCF: data_out = 8'hCE;
                    16'hFFD0: data_out = 8'hCF;
                    16'hFFD1: data_out = 8'hD0;
                    16'hFFD2: data_out = 8'hD1;
                    16'hFFD3: data_out = 8'hD2;
                    16'hFFD4: data_out = 8'hD3;
                    16'hFFD5: data_out = 8'hD4;
                    16'hFFD6: data_out = 8'hD5;
                    16'hFFD7: data_out = 8'hD6;
                    16'hFFD8: data_out = 8'hD7;
                    16'hFFD9: data_out = 8'hD8;
                    16'hFFDA: data_out = 8'hD9;
                    16'hFFDB: data_out = 8'hDA;
                    16'hFFDC: data_out = 8'hDB;
                    16'hFFDD: data_out = 8'hDC;
                    16'hFFDE: data_out = 8'hDD;
                    16'hFFDF: data_out = 8'hDE;
                    16'hFFE0: data_out = 8'hDF;
                    16'hFFE1: data_out = 8'hE0;
                    16'hFFE2: data_out = 8'hE1;
                    16'hFFE3: data_out = 8'hE2;
                    16'hFFE4: data_out = 8'hE3;
                    16'hFFE5: data_out = 8'hE4;
                    16'hFFE6: data_out = 8'hE5;
                    16'hFFE7: data_out = 8'hE6;
                    16'hFFE8: data_out = 8'hE7;
                    16'hFFE9: data_out = 8'hE8;
                    16'hFFEA: data_out = 8'hE9;
                    16'hFFEB: data_out = 8'hEA;
                    16'hFFEC: data_out = 8'hEB;
                    16'hFFED: data_out = 8'hEC;
                    16'hFFEE: data_out = 8'hED;
                    16'hFFEF: data_out = 8'hEE;
                    16'hFFF0: data_out = 8'hEF;
                    16'hFFF1: data_out = 8'hF0;
                    16'hFFF2: data_out = 8'hF1;
                    16'hFFF3: data_out = 8'hF2;
                    16'hFFF4: data_out = 8'hF3;
                    16'hFFF5: data_out = 8'hF4;
                    16'hFFF6: data_out = 8'hF5;
                    16'hFFF7: data_out = 8'hF6;
                    16'hFFF8: data_out = 8'hF7;
                    16'hFFF9: data_out = 8'hF8;
                    16'hFFFA: data_out = 8'hF9;
                    16'hFFFB: data_out = 8'hFA;
                    16'hFFFC: data_out = 8'hFB;
                    16'hFFFD: data_out = 8'hFC;
                    16'hFFFE: data_out = 8'hFD;
                    16'hFFFF: data_out = 8'hFE;
                    default: data_out = 8'h00;
                endcase
            end
        end
    endgenerate

    always_ff @( posedge clk ) 
    begin
        adder_out <= data_out;
    end

endmodule