module fwft #( //First Word Fall Through
    parameter  DATA_WIDTH = 32,
    parameter  ADDR_WIDTH = 4,
    localparam OUT_WIDTH  = DATA_WIDTH >> 1
)(
    input  logic                  clk,
    input  logic                  arst_n,

    // Write Interface
    input  logic                  wr,
    input  logic [DATA_WIDTH-1:0] wr_data,
    output logic                  full,

    // Read Interface
    input  logic                  rd,
    output logic [OUT_WIDTH-1:0]  rd_data,
    output logic                  empty
);

    logic [ADDR_WIDTH-1:0] ctrl_wr_addr;
    logic [ADDR_WIDTH-1:0] ctrl_rd_addr;
    logic                  byte_rd;
    
    logic [DATA_WIDTH-1:0] rf_rd_data;

    logic                  ctrl_wr_en;
    logic                  ctrl_full;

    assign ctrl_wr_en = wr & !ctrl_full;
    assign full       = ctrl_full;
    assign rd_data    = byte_rd ? rf_rd_data[OUT_WIDTH +: OUT_WIDTH] : rf_rd_data[OUT_WIDTH-1 : 0];

    fifo_ctrl #(
        .ADDR_WIDTH( ADDR_WIDTH )
    ) u_fifo_ctrl (
        .clk    ( clk          ),
        .arst_n ( arst_n       ),
        .wr_en  ( wr           ),
        .wr_addr( ctrl_wr_addr ),
        .full   ( ctrl_full    ),
        .rd_en  ( rd           ),
        .byte_rd( byte_rd      ),
        .rd_addr( ctrl_rd_addr ),
        .empty  ( empty        )
    );

    register_file #(
        .DATA_WIDTH( DATA_WIDTH ),
        .ADDR_WIDTH( ADDR_WIDTH )
    ) u_reg_file (
        .clk    ( clk          ),
        .arst_n ( arst_n       ),
        .wr_en  ( ctrl_wr_en   ),
        .wr_data( wr_data      ),
        .wr_addr( ctrl_wr_addr ),
        .rd_addr( ctrl_rd_addr ),
        .rd_data( rf_rd_data   )
    );
    
endmodule